
GS1 i LUTs

constant lut_gs_1 : vector_of_std_logic_vector16(0 to 63) := 
  ("0000000010001011",
   "0010101011011001",
   "0010001101101001",
   "1110000010101001",
   "1101110010100010",
   "1110000000100100",
   "1101111101010101",
   "1101111011000100",
   "1101110001111110",
   "0001111001000001",
   "1110001110000001",
   "0010000000001100",
   "0001110101001110",
   "1101111011010000",
   "0010010111101100",
   "0010000111000001",
   "0010000010101011",
   "0010000000100101",
   "0001111000111111",
   "1110000100111010",
   "0010000111000001",
   "1101110110101110",
   "1110001011010111",
   "0001110110010111",
   "0001101000111010",
   "0010000010101011",
   "0001110100101001",
   "1101110100000100",
   "0001101001010011",
   "1101100110001101",
   "0010001011001101",
   "0010010010111101",
   "0010010000101100",
   "0001111101010111",
   "1101110001011011",
   "1101100011111110",
   "0001111011101011",
   "0010000011110100",
   "1101101101000011",
   "0010000100110000",
   "0001101000111010",
   "0001101010011011",
   "1101110110101110",
   "0010010010111101",
   "0010000000000001",
   "1101110110101110",
   "0010000110011100",
   "1110000100001011",
   "0001111000011100",
   "1110000001100000",
   "1110011100000001",
   "0010010010011000",
   "0010010010001101",
   "1101011010110111",
   "0010000110011110",
   "0010000100010111",
   "1101100100111010",
   "1101111111100110",
   "1101100010010000",
   "1110001001000110",
   "0010011111110101",
   "1110011011011101",
   "1110010110101101",
   "0010001110100111");



constant lut_gs_2 : vector_of_std_logic_vector16(0 to 63) := 
  ("0000000001110111",
   "0010011101110011",
   "0001101010101101",
   "1110010110111011",
   "1101110010011000",
   "1110011111001100",
   "1110001001001011",
   "1110011100111101",
   "1101010000100101",
   "0001001101001110",
   "1110001001101101",
   "0001111100010000",
   "0010001100010100",
   "1110011100000001",
   "0010000001101110",
   "0001110110110101",
   "0001010000001100",
   "0001101101110100",
   "0001110011101001",
   "1101101110100001",
   "0010100111010011",
   "1110011001001111",
   "1110000001100101",
   "0001001001000010",
   "0001111010001011",
   "0010010110011011",
   "0001110011101001",
   "1101011111000000",
   "0001101011101110",
   "1101111000001010",
   "0010001011001100",
   "0010101001001000",
   "0001110101111000",
   "0010001100100111",
   "1101101000110011",
   "1101111110010010",
   "0010011111011000",
   "0001101111000000",
   "1101001111110101",
   "0010011111011100",
   "0001110110011100",
   "0010001010010100",
   "1101011101100101",
   "0001110100101110",
   "0010100011000111",
   "1110010101010011",
   "0010011001100111",
   "1110000011110000",
   "0001010001110101",
   "1101111111010110",
   "1110010011100001",
   "0001110011111110",
   "0010001001111101",
   "1101011000010100",
   "0001110011001100",
   "0010101100011101",
   "1101110011010001",
   "1110011100000001",
   "1101110100011111",
   "1101111000000101",
   "0010000010000001",
   "1110001001100100",
   "1110011000001110",
   "0001110000110011");



constant lut_gs_3 : vector_of_std_logic_vector16(0 to 63) := 
  ("0000000001000011",
   "0001111000110101",
   "0001000010000100",
   "1110101101100101",
   "1110000101010100",
   "1110111110110011",
   "1110011110101011",
   "1111000111101001",
   "1100111101001000",
   "0000011101110000",
   "1101111110001100",
   "0001111011000100",
   "0010100001111011",
   "1110111110101111",
   "0001011101111111",
   "0001100001010101",
   "0000011000010011",
   "0001100000100000",
   "0001110101000011",
   "1101011111010101",
   "0010111011010010",
   "1111000101100010",
   "1101110110100110",
   "0000011101110000",
   "0010001101100001",
   "0010100000011101",
   "0001110101000011",
   "1101010111001011",
   "0001110010111101",
   "1110011101111111",
   "0001111001111011",
   "0010110000011011",
   "0001010100010010",
   "0010011001001010",
   "1101100001011011",
   "1110100010000001",
   "0010111001001011",
   "0001010000111101",
   "1100111101010101",
   "0010110101000100",
   "0010001011011010",
   "0010100110000111",
   "1101001100001111",
   "0001001110111000",
   "0010111011010010",
   "1110111101111100",
   "0010101000010001",
   "1110000100111100",
   "0000101100110111",
   "1101111111011100",
   "1110000101100000",
   "0001001111000101",
   "0001110100011110",
   "1101101110110100",
   "0001010000111101",
   "0011001000010101",
   "1110010010010101",
   "1110111110101111",
   "1110010111110001",
   "1101100011100101",
   "0001010101001110",
   "1101110100100110",
   "1110010100101001",
   "0001000111010001");



constant lut_gs_4 : vector_of_std_logic_vector16(0 to 63) := 
  ("1111111111110110",
   "0001000010000010",
   "0000010100101011",
   "1111001000011111",
   "1110100111000011",
   "1111100000011110",
   "1110111011001001",
   "1111110101101101",
   "1100110101110101",
   "1111101111111111",
   "1101110000000100",
   "0001111010011001",
   "0010110101010001",
   "1111100011101100",
   "0000110001011001",
   "0001000100110111",
   "1111100001110000",
   "0001010111111010",
   "0001111010001000",
   "1101010101111010",
   "0011000100011011",
   "1111110110000001",
   "1101101010010100",
   "1111110100111010",
   "0010100001110110",
   "0010100011011101",
   "0001111010001000",
   "1101011001001011",
   "0001111111011000",
   "1111010000011111",
   "0001011011010110",
   "0010101100100101",
   "0000101011111101",
   "0010100000110011",
   "1101011110001110",
   "1111001110100111",
   "0011001001101011",
   "0000101010101001",
   "1100110111100010",
   "0011000010011101",
   "0010100010001010",
   "0010111101010000",
   "1101000100111000",
   "0000100010010101",
   "0011001001010111",
   "1111101011010101",
   "0010101111110111",
   "1110000101100111",
   "0000001000111001",
   "1101111111100011",
   "1101110010101110",
   "0000100100000011",
   "0001010010000011",
   "1110011000111000",
   "0000100101101110",
   "0011011000011001",
   "1111000000010010",
   "1111100011101100",
   "1111001001100101",
   "1101010000110100",
   "0000011100111011",
   "1101011101110110",
   "1110001011010100",
   "0000010111101001");



constant lut_gs_5 : vector_of_std_logic_vector16(0 to 63) := 
  ("1111111110011100",
   "0000000001100100",
   "1111100110011100",
   "1111100111001001",
   "1111010011110101",
   "0000000011001000",
   "1111011101011011",
   "0000100011010010",
   "1100111001110110",
   "1111000110111111",
   "1101100010100011",
   "0001111010001011",
   "0011000011001001",
   "0000001000111001",
   "0000000000000000",
   "0000100010100101",
   "1110110001010000",
   "0001010100111101",
   "0010000001001000",
   "1101010010101101",
   "0011000011000010",
   "0000100110011010",
   "1101011111011011",
   "1111010000101101",
   "0010110011001100",
   "0010100000100101",
   "0010000001001000",
   "1101100010100011",
   "0010001101111110",
   "0000001000111001",
   "0000110010011011",
   "0010100000100101",
   "0000000000000000",
   "0010100011101101",
   "1101011111011011",
   "0000000000000000",
   "0011001111111000",
   "0000000000000000",
   "1100111100110111",
   "0011000110111110",
   "0010110110010100",
   "0011001100110000",
   "1101000110100100",
   "1111110011010001",
   "0011001100110000",
   "0000011001100100",
   "0010110000011011",
   "1110000101110101",
   "1111100111001001",
   "1101111111100101",
   "1101011111011011",
   "1111110110010010",
   "0000100110011010",
   "1111010000101101",
   "1111110110010010",
   "0011011011111001",
   "1111110111000111",
   "0000001000111001",
   "0000000011001000",
   "1101000011000111",
   "1111100000100011",
   "1101001001101100",
   "1101111110111000",
   "1111100110011100");



constant lut_gs_6 : vector_of_std_logic_vector16(0 to 63) := 
  ("1111111101001000",
   "1111000001000000",
   "1110111011100111",
   "0000001000111001",
   "0000000110110001",
   "0000100101100111",
   "0000000011111110",
   "0001001100010011",
   "1101000111010111",
   "1110100101011111",
   "1101011001001011",
   "0001111010011001",
   "0011001000011110",
   "0000101100100001",
   "1111001110100111",
   "1111111100000010",
   "1110001011001010",
   "0001010111111010",
   "0010000111111001",
   "1101010101111010",
   "0010111000010101",
   "0001010010000011",
   "1101011000110111",
   "1110110010110101",
   "0010111101011110",
   "0010011001011000",
   "0010000111111001",
   "1101110000000100",
   "0010011010111111",
   "0000111111101110",
   "0000000011000000",
   "0010010000010000",
   "1111010100000011",
   "0010100010000111",
   "1101100100111101",
   "0000110001011001",
   "0011001011011011",
   "1111010101010111",
   "1101001010101111",
   "0011000010011101",
   "0011000011001110",
   "0011010001110001",
   "1101001111101011",
   "1111000110010011",
   "0011000101101011",
   "0001000100011001",
   "0010101010011011",
   "1110000101100111",
   "1111001000011111",
   "1101111111100011",
   "1101010000011100",
   "1111001001101100",
   "1111110110000001",
   "0000001110110111",
   "1111001000000000",
   "0011010010111110",
   "0000101111100001",
   "0000101100100001",
   "0000111100100000",
   "1100111101100111",
   "1110101000010000",
   "1100111100110010",
   "1101110010101011",
   "1110111000101001");



constant lut_gs_7 : vector_of_std_logic_vector16(0 to 63) := 
  ("1111111100001101",
   "1110001001111011",
   "1110011000010101",
   "0000101100110111",
   "0000111010100001",
   "0001000110101101",
   "0000101100110111",
   "0001101100111000",
   "1101011100000000",
   "1110001101101100",
   "1101010111001011",
   "0001111011000100",
   "0011000010101011",
   "0001001100111011",
   "1110100010000001",
   "1111010011001001",
   "1101110011000100",
   "0001100000100000",
   "0010001100000111",
   "1101011111010101",
   "0010100110000111",
   "0001110100011110",
   "1101011001010010",
   "1110011100100110",
   "0010111101001011",
   "0010001111101011",
   "0010001100000111",
   "1101111110001100",
   "0010100010100111",
   "0001101101101011",
   "1111010001010000",
   "0001111111101101",
   "1110101011101110",
   "0010011100011110",
   "1101101110011101",
   "0001011101111111",
   "0010111100100111",
   "1110101111000011",
   "1101011110000101",
   "0010110101000100",
   "0011000100110010",
   "0011001010001100",
   "1101011110000101",
   "1110011111111100",
   "0010110101000001",
   "0001100111101011",
   "0010011110100100",
   "1110000100111100",
   "1110101101100101",
   "1101111111011100",
   "1101001010011000",
   "1110100010000001",
   "1111000101100010",
   "0001001011100010",
   "1110100000001001",
   "0010111110101000",
   "0001100010000001",
   "0001001100111011",
   "0001101101101111",
   "1101000010110101",
   "1101111011110101",
   "1100111011001110",
   "1101101010001100",
   "1110010011001000");



constant lut_gs_8 : vector_of_std_logic_vector16(0 to 63) := 
  ("1111111011111100",
   "1101100100011010",
   "1110000000000100",
   "0001010001110101",
   "0001101001111100",
   "0001100101001110",
   "0001010110000010",
   "0010000001110101",
   "1101110101001110",
   "1110000001001001",
   "1101011111000000",
   "0001111100010000",
   "0010110000001011",
   "0001101000111000",
   "1101111110010010",
   "1110101001111110",
   "1101101011010101",
   "0001101101110100",
   "0010001011101001",
   "1101101110100001",
   "0010001110100001",
   "0010001001111101",
   "1101100010101111",
   "1110001110111001",
   "0010101111111110",
   "0010000101010001",
   "0010001011101001",
   "1110001001101101",
   "0010100001100010",
   "0010001100101111",
   "1110100001010011",
   "0001110010100100",
   "1110001010001000",
   "0010010011011111",
   "1101111011100001",
   "0010000001101110",
   "0010100100011001",
   "1110010001000000",
   "1101110011101100",
   "0010011111011100",
   "0010111000000110",
   "0010110101000011",
   "1101101111011111",
   "1110000100000000",
   "0010011100010001",
   "0001111111111100",
   "0010001101110000",
   "1110000011110000",
   "1110010110111011",
   "1101111111010110",
   "1101010000110011",
   "1110000010011110",
   "1110011001001111",
   "0001111111100111",
   "1110000011010000",
   "0010100000100111",
   "0010000111110110",
   "0001101000111000",
   "0010001111111010",
   "1101010100001110",
   "1101100001100101",
   "1101000111111010",
   "1101101000100000",
   "1101111001111111");



constant lut_gs_9 : vector_of_std_logic_vector16(0 to 63) := 
  ("1111111010010101",
   "1101010011110001",
   "1101110111011101",
   "0001111000011100",
   "0010001110100111",
   "0010000010000110",
   "0001111111011100",
   "0010001011001101",
   "1110010010111011",
   "1101111110011101",
   "1101101111101101",
   "0001111011110101",
   "0010001110100111",
   "0001111101010111",
   "1101100011111110",
   "1110000100111010",
   "1101110110111000",
   "0010000000100101",
   "0010000010101011",
   "1110000000100100",
   "0001110101110010",
   "0010001101110111",
   "1101111000011010",
   "1110001000001000",
   "0010010111010011",
   "0001111101111010",
   "0010000111000001",
   "1110010010010111",
   "0010010011010110",
   "0010011011000110",
   "1101110100101000",
   "0001101001010011",
   "1101110011101011",
   "0010001010001111",
   "1110001101111111",
   "0010010111101100",
   "0010000110011100",
   "1110000000100010",
   "1110001010110010",
   "0010000000011010",
   "0010011110010011",
   "0010010101000010",
   "1101111111011011",
   "1101110011000111",
   "0001111111011100",
   "0010001100111001",
   "0001111011000110",
   "1110000100001011",
   "1110000110111111",
   "1101111101001010",
   "1101100011011001",
   "1101101111010100",
   "1101110110101110",
   "0010100111111110",
   "1101110010100010",
   "0001111101010111",
   "0010011001110011",
   "0010000001101101",
   "0010100000011010",
   "1101110100000100",
   "1101011111100110",
   "1101100001101101",
   "1101101101101000",
   "1101110010001001");



constant lut_gs_10 : vector_of_std_logic_vector16(0 to 63) := 
  ("1111111100000011",
   "1101011110100111",
   "1101111100111101",
   "0010011000000100",
   "0010101100010000",
   "0010011001100111",
   "0010100000001101",
   "0010000101100011",
   "1110101100101111",
   "1110001000001101",
   "1110001111101011",
   "0001111100011101",
   "0001100110000001",
   "0010001100100111",
   "1101011010110000",
   "1101100011100010",
   "1110001110000010",
   "0010010100001111",
   "0001110110110101",
   "1110011011010000",
   "0001010111000000",
   "0010000110000001",
   "1110010011011010",
   "1110001011001011",
   "0001101101101011",
   "0001110100001100",
   "0001111010100100",
   "1110010100010010",
   "0001111110000000",
   "0010010000101011",
   "1101010100110001",
   "0001101011101110",
   "1101100010101011",
   "0001111111010010",
   "1110011111000011",
   "0010100001100010",
   "0001011110001010",
   "1101111001000101",
   "1110011010010101",
   "0001100000000011",
   "0001110001110111",
   "0001100101100111",
   "1110001110011110",
   "1101110101010010",
   "0001011001111110",
   "0010000110110010",
   "0001100100110000",
   "1110000011100011",
   "1101110111010101",
   "1101111011101000",
   "1110000100100101",
   "1101100110100111",
   "1101011101100101",
   "0010111011000100",
   "1101110010011000",
   "0001010100111001",
   "0010011011110101",
   "0010010000010110",
   "0010011010011111",
   "1110011110001100",
   "1101110100000010",
   "1110001110001001",
   "1110000001010000",
   "1101110110000011");



constant lut_gs_11 : vector_of_std_logic_vector16(0 to 63) := 
  ("1111111110111101",
   "1110000001010001",
   "1110001101101100",
   "0010110101000001",
   "0010111011000101",
   "0010101000010001",
   "0010111100100111",
   "0001101110111110",
   "1111001000001101",
   "1110011111111100",
   "1110110110101000",
   "0010000000100100",
   "0000110010111011",
   "0010011001001010",
   "1101011011010010",
   "1101000101011111",
   "1110110100011111",
   "0010100100000001",
   "0001100001010101",
   "1110110111001100",
   "0000111001111010",
   "0001101100111000",
   "1110111000101111",
   "1110011010011111",
   "0000111100101000",
   "0001101111010110",
   "0001100011011011",
   "1110001101000011",
   "0001011011111000",
   "0001110101010001",
   "1100111101001000",
   "0001110010111101",
   "1101011101011001",
   "0001110001100000",
   "1110110101001100",
   "0010100010100111",
   "0000110100011101",
   "1110000001111110",
   "1110100111000111",
   "0000111001101011",
   "0000111100101000",
   "0000110000111010",
   "1110011101011010",
   "1110000011111111",
   "0000110100011101",
   "0001110100011011",
   "0001001000110100",
   "1101111111011100",
   "1101101110011101",
   "1101111101010110",
   "1110110100011110",
   "1101100100111111",
   "1101001100001111",
   "0010111111010101",
   "1110000101010100",
   "0000100111011101",
   "0010000111011111",
   "0010011011010000",
   "0001111100100101",
   "1111001101000101",
   "1110011001111000",
   "1111000011011000",
   "1110011100100101",
   "1110001011100010");



constant lut_gs_12 : vector_of_std_logic_vector16(0 to 63) := 
  ("0000000010101000",
   "1110110110011110",
   "1110101010011010",
   "0011001010100110",
   "0010111101110010",
   "0010101111110111",
   "0011010000010111",
   "0001001011111110",
   "1111100010110100",
   "1111000001011000",
   "1111100011101111",
   "0010000101011001",
   "1111111100000101",
   "0010100000110011",
   "1101100101010101",
   "1100101111010101",
   "1111100011100101",
   "0010110000000000",
   "0001000100110111",
   "1111010101110010",
   "0000011100111000",
   "0001000111010111",
   "1111100011011011",
   "1110110011001001",
   "0000000110011101",
   "0001101101011010",
   "0001000100100011",
   "1110000000101000",
   "0000110001101101",
   "0001001010011010",
   "1100110000111001",
   "0001111111011000",
   "1101100000000101",
   "0001100100111100",
   "1111001110001111",
   "0010011010111111",
   "0000001001101110",
   "1110011000100000",
   "1110101101110110",
   "0000010001101000",
   "0000000001100001",
   "1111111001011110",
   "1110101000011010",
   "1110100000000011",
   "0000001110101010",
   "0001010101010001",
   "0000101010001110",
   "1101111010100111",
   "1101101001111001",
   "1101111111110111",
   "1111101100001101",
   "1101101010110001",
   "1101000100111000",
   "0010110101000000",
   "1110100111000011",
   "1111111010010110",
   "0001100001101100",
   "0010100000011111",
   "0001001101000100",
   "1111111110111111",
   "1111001110001100",
   "1111111110011111",
   "1111000000011001",
   "1110101101111101");



constant lut_gs_13 : vector_of_std_logic_vector16(0 to 63) := 
  ("0000000110011011",
   "1111110110010010",
   "1111010000101101",
   "0011010110011101",
   "0010110110010100",
   "0010110000011011",
   "0011011001100101",
   "0000100000001010",
   "1111111100111000",
   "1111101001100100",
   "0000010010111111",
   "0010001010001000",
   "1111000110111111",
   "0010100011101101",
   "1101110101001010",
   "1100100011010011",
   "0000010101101111",
   "0010110110010100",
   "0000100010100101",
   "1111110110010010",
   "0000000000000000",
   "0000011001100100",
   "0000001111110111",
   "1111010011110101",
   "1111010000101101",
   "0001101110001001",
   "0000011111011101",
   "1101110010000010",
   "0000000011001000",
   "0000010101101111",
   "1100110000001000",
   "0010001101111110",
   "1101101000010101",
   "0001011011100010",
   "1111101010010001",
   "0010001101111110",
   "1111100000100011",
   "1110111010111110",
   "1110101110001011",
   "1111101010010001",
   "1111000110111111",
   "1111000100101011",
   "1110101110001011",
   "1111000110111111",
   "1111101010010001",
   "0000101100001011",
   "0000001001101110",
   "1101110101111000",
   "1101101001001001",
   "1110000010101101",
   "0000100101100110",
   "1101110101001010",
   "1101000110100100",
   "0010100000100101",
   "1111010011110101",
   "1111010000101101",
   "0000101111010011",
   "0010100000100101",
   "0000010010100111",
   "0000101111010011",
   "0000001001101110",
   "0000111001000001",
   "1111101010010001",
   "1111011001100110");



constant lut_gs_14 : vector_of_std_logic_vector16(0 to 63) := 
  ("0000001001100011",
   "0000110111010000",
   "1111111101010101",
   "0011010110101101",
   "0010100111100110",
   "0010101010011011",
   "0011010111000001",
   "1111101111111100",
   "0000010111001000",
   "0000010100111111",
   "0000111111110001",
   "0010001101110011",
   "1110011001011000",
   "0010100010000111",
   "1110000110011001",
   "1100100011001111",
   "0001000100111110",
   "0010110101011000",
   "1111111100000010",
   "0000010111111100",
   "1111100011001000",
   "1111101000010111",
   "0000111010000001",
   "1111111010101011",
   "1110100001010011",
   "0001110001000110",
   "1111110110010010",
   "1101100101000001",
   "1111010100011000",
   "1111011110001001",
   "1100111010000001",
   "0010011010111111",
   "1101110011010010",
   "0001010111000110",
   "0000001001001110",
   "0001111111011000",
   "1110111011011101",
   "1111100110101100",
   "1110101000011010",
   "1111000101110101",
   "1110010011111101",
   "1110011000000000",
   "1110101101110110",
   "1111110101011011",
   "1111001000110011",
   "1111111100111011",
   "1111101000000100",
   "1101110010001101",
   "1101101011100100",
   "1110000101010011",
   "0001011001110010",
   "1110000000111101",
   "1101001111101011",
   "0010000111110110",
   "0000000110110001",
   "1110101101011001",
   "1111110110100101",
   "0010011100010110",
   "1111010101011010",
   "0001011001010001",
   "0001000100000110",
   "0001101100000011",
   "0000010111000100",
   "0000001001111111");



constant lut_gs_15 : vector_of_std_logic_vector16(0 to 63) := 
  ("0000001011010000",
   "0001101111110101",
   "0000101100101010",
   "0011001010001100",
   "0010010101000111",
   "0010011110100100",
   "0011001000000101",
   "1111000000000011",
   "0000110010010011",
   "0000111111111101",
   "0001100101100100",
   "0010001111011110",
   "1101111000100001",
   "0010011100011110",
   "1110010100101001",
   "1100110000010100",
   "0001101011100101",
   "0010101100001011",
   "1111010011001001",
   "0000111001111010",
   "1111000110000110",
   "1110111000101111",
   "0001011101111110",
   "0000100101010110",
   "1101111101101110",
   "0001110101100111",
   "1111001011100011",
   "1101011101011001",
   "1110101001101000",
   "1110101010110010",
   "1101001101000101",
   "0010100010100111",
   "1101111110001001",
   "0001011000111001",
   "0000101010110001",
   "0001110010111101",
   "1110011100100101",
   "0000011000010011",
   "1110011101011010",
   "1110100110010010",
   "1101101110110100",
   "1101111000010001",
   "1110100111000111",
   "0000100111011101",
   "1110101011011111",
   "1111001011110000",
   "1111000110000110",
   "1101110000100010",
   "1101110000010101",
   "1110000111000011",
   "0010000010010010",
   "1110001010111101",
   "1101011110000101",
   "0001110000110011",
   "0000111010100001",
   "1110010010111001",
   "1110111110001011",
   "0010010100111000",
   "1110011101111111",
   "0001111000100101",
   "0001110101000010",
   "0010010001001100",
   "0001000011010111",
   "0000111010011110");



constant lut_gs_16 : vector_of_std_logic_vector16(0 to 63) := 
  ("0000001010111100",
   "0010010111110101",
   "0001011010111110",
   "0010110000110111",
   "0010000010010011",
   "0010001101110000",
   "0010101101001000",
   "1110010100110101",
   "0001001110110111",
   "0001100110111110",
   "0010000000011010",
   "0010001110011010",
   "1101101000010111",
   "0010010011011111",
   "1110011100011010",
   "1101001010110000",
   "0010000100110100",
   "0010011010010011",
   "1110101001111110",
   "0001011011001100",
   "1110101001000000",
   "1110001111001101",
   "0001111000010001",
   "0001010001001010",
   "1101101010010000",
   "0001111011000010",
   "1110100001110110",
   "1101011110011110",
   "1110000110011010",
   "1110000010001011",
   "1101100111011110",
   "0010100001100010",
   "1110000110100010",
   "0001100001011111",
   "0001001110000111",
   "0001101011101110",
   "1110000101011100",
   "0001001100000000",
   "1110001110011110",
   "1110001101000110",
   "1101011100100000",
   "1101101001000010",
   "1110011010010101",
   "0001011001000101",
   "1110010011001100",
   "1110011100111001",
   "1110100100110100",
   "1101110001100110",
   "1101110110100011",
   "1110000111011110",
   "0010011001111100",
   "1110010000100011",
   "1101101111011111",
   "0001100000101000",
   "0001101001111100",
   "1110000011000010",
   "1110001100001111",
   "0010001011010111",
   "1101110011111101",
   "0010001001111001",
   "0010010101100010",
   "0010100011100000",
   "0001101011111010",
   "0001100110110001");



constant lut_gs_17 : vector_of_std_logic_vector16(0 to 63) := 
  ("0000001010100000",
   "0010100111011010",
   "0010000111000001",
   "0010001001101011",
   "0001110100010000",
   "0001111011000110",
   "0010001001101011",
   "1101101111101101",
   "0001101010011011",
   "0010001001010010",
   "0010001011001101",
   "0010001000001010",
   "1101101101001110",
   "0010000101111001",
   "1110011001010111",
   "1101101111010100",
   "0010001011011001",
   "0001111101111100",
   "1110000000100100",
   "0001111100110010",
   "1110001110100100",
   "1101110001011001",
   "0010000100001101",
   "0001111001000001",
   "1101101011100010",
   "0001111110011111",
   "1101111001100100",
   "1101101000010100",
   "1101101010111110",
   "1101101011100010",
   "1110001001010000",
   "0010010011010110",
   "1110001101000011",
   "0001110010100100",
   "0001110100000110",
   "0001101101101001",
   "1101111000111111",
   "0001111011101011",
   "1101111111011011",
   "1101111000111111",
   "1101100001110111",
   "1101101001110101",
   "1110000110011100",
   "0010001000101110",
   "1110000010101001",
   "1101110110010101",
   "1110000111100100",
   "1101110011100000",
   "1101111111011011",
   "1110001000100001",
   "0010011011011111",
   "1110010010010111",
   "1101111111011011",
   "0001011100111110",
   "0010010010111101",
   "1101111100110001",
   "1101100111101111",
   "0001111110111000",
   "1101011111001101",
   "0010001101011110",
   "0010100011000100",
   "0010100010011111",
   "0010001011110001",
   "0010001001010010");



constant lut_gs_18 : vector_of_std_logic_vector16(0 to 63) := 
  ("0000000101011100",
   "0010011110111001",
   "0010101011001111",
   "0001011001110000",
   "0001100110011100",
   "0001100100110000",
   "0001011101011110",
   "1101010101101010",
   "0010000110100110",
   "0010100010001110",
   "0010001011001100",
   "0010000011101000",
   "1110000000010010",
   "0001111011100100",
   "1110001101111010",
   "1110011110010101",
   "0010000100110100",
   "0001011110110110",
   "1101011111110011",
   "0010010110101001",
   "1101110101001110",
   "1101011010100111",
   "0010000110111111",
   "0010100000100111",
   "1101111111000100",
   "0010000010000101",
   "1101011011100111",
   "1101111110010010",
   "1101011110111100",
   "1101100111001001",
   "1110101001110001",
   "0001111110000000",
   "1110001010011110",
   "0010000111111011",
   "0010011000000100",
   "0001110110010011",
   "1101110100010111",
   "0010101010001010",
   "1101101111011111",
   "1101101100101100",
   "1101111100000110",
   "1110000000111101",
   "1101101111111101",
   "0010101100011101",
   "1101110111010101",
   "1101010100010011",
   "1101101101000101",
   "1101111000101010",
   "1110000111011010",
   "1110000011100011",
   "0010001001000101",
   "1110001101011100",
   "1110001110011110",
   "0001100100010110",
   "0010101111111110",
   "1110000110111110",
   "1101001100110111",
   "0001110111010111",
   "1101011100000010",
   "0010000000011110",
   "0010011001010001",
   "0010000111101001",
   "0010100011101001",
   "0010100010011011");



constant lut_gs_19 : vector_of_std_logic_vector16(0 to 63) := 
  ("1111111110010101",
   "0010000010000101",
   "0011000010111000",
   "0000100111001101",
   "0001100000011100",
   "0001001000110100",
   "0000101001010100",
   "1101001010001001",
   "0010100100000000",
   "0010101110010001",
   "0001111001111011",
   "0001111011000111",
   "1110100101100101",
   "0001101111011010",
   "1101111110001100",
   "1111010110101100",
   "0001101011100101",
   "0000111000010111",
   "1101000011011001",
   "0010101101101101",
   "1101011100000000",
   "1101010001101011",
   "0001111001111011",
   "0010111110101000",
   "1110100000001001",
   "0010000111110111",
   "1101000011011001",
   "1110100010000001",
   "1101011011010010",
   "1101110011000100",
   "1111001101101001",
   "0001011011111000",
   "1110000101101111",
   "0010011100011011",
   "0010110101000001",
   "0010000001110100",
   "1101110011111001",
   "0011001101100010",
   "1101011110000101",
   "1101101010001100",
   "1110100101100101",
   "1110100101010110",
   "1101011011111111",
   "0011001000010101",
   "1101101110011101",
   "1100111111001110",
   "1101010100011001",
   "1110000010110010",
   "1110001011001010",
   "1101111111011100",
   "0001100111011110",
   "1110000000010011",
   "1110011101011010",
   "0001110010111010",
   "0010111101001011",
   "1110011010011111",
   "1101000010110001",
   "0001101111011010",
   "1101110000111010",
   "0001100001111110",
   "0001110111001001",
   "0001011100100001",
   "0010110101000100",
   "0010110011110001");



constant lut_gs_20 : vector_of_std_logic_vector16(0 to 63) := 
  ("1111110110010001",
   "0001010011001001",
   "0011001111000111",
   "1111110100000010",
   "0001100000000100",
   "0000101010001110",
   "1111110011101110",
   "1101001010001000",
   "0010111101100101",
   "0010110000001000",
   "0001011011010110",
   "0001110010001111",
   "1111010110001111",
   "0001100101010000",
   "1101101011001001",
   "0000010001001110",
   "0001000100111110",
   "0000001111001111",
   "1100101111101001",
   "0010111110000101",
   "1101000111010111",
   "1101010011000110",
   "0001100000010001",
   "0011010010111110",
   "1111001100111100",
   "0010001100111111",
   "1100110100100101",
   "1111001110100111",
   "1101100000011001",
   "1110010000000110",
   "1111110001000010",
   "0000110001101101",
   "1101111101111110",
   "0010101111001100",
   "0011001010100110",
   "0010001111111100",
   "1101111000000111",
   "0011100101001111",
   "1101001111101011",
   "1101101101101111",
   "1111011011001010",
   "1111010100110110",
   "1101001011000100",
   "0011011000011001",
   "1101101001111001",
   "1100110101100000",
   "1101000001100111",
   "1110001110000110",
   "1110001100100001",
   "1101111010100111",
   "0000111000110100",
   "1101101111110000",
   "1110101000011010",
   "0010000111100001",
   "0010111101011110",
   "1110111000000101",
   "1101000101110000",
   "0001101010001100",
   "1110011000100100",
   "0000110111101011",
   "0001000011110001",
   "0000100100100001",
   "0010111101100001",
   "0010111011001000");



constant lut_gs_21 : vector_of_std_logic_vector16(0 to 63) := 
  ("1111101110101110",
   "0000011000110111",
   "0011001111111000",
   "1111000100101011",
   "0001100100011100",
   "0000001001101110",
   "1111000001100011",
   "1101010011011010",
   "0011001111111000",
   "0010101001011110",
   "0000110010011011",
   "0001101010101100",
   "0000001100000001",
   "0001011110101010",
   "1101011000110110",
   "0001001000001010",
   "0000010101101111",
   "1111100110011100",
   "1100100110011011",
   "0011000110001010",
   "1100111001110110",
   "1101011100010011",
   "0000111100001001",
   "0011011011111001",
   "0000000000000000",
   "0010010000101110",
   "1100110000001000",
   "0000000000000000",
   "1101101011011101",
   "1110111010111110",
   "0000010010100111",
   "0000000011001000",
   "1101110101001010",
   "0010111100111001",
   "0011010110011101",
   "0010011101011101",
   "1101111110111000",
   "0011101111010100",
   "1101000110100100",
   "1101110101001010",
   "0000010101101111",
   "0000001001101110",
   "1100111111111111",
   "0011011011111001",
   "1101101001001001",
   "1100110110101110",
   "1100110110101110",
   "1110011000011100",
   "1110001011100111",
   "1101110101111000",
   "0000000011001000",
   "1101011111011011",
   "1110101110001011",
   "0010011101011101",
   "0010110011001100",
   "1111011101100010",
   "1101010010100110",
   "0001101000011000",
   "1111001101100101",
   "0000000110100110",
   "0000000110100110",
   "1111100111001001",
   "0010111101010001",
   "0010111001011100");



constant lut_gs_22 : vector_of_std_logic_vector16(0 to 63) := 
  ("1111101001010011",
   "1111011011011111",
   "0011000101111111",
   "1110011101011100",
   "0001101100001010",
   "1111101000000100",
   "1110010111101100",
   "1101100010110001",
   "0011010111100001",
   "0010011100111010",
   "0000000011000000",
   "0001100110001001",
   "0001000000000010",
   "0001011100110110",
   "1101001011110101",
   "0001110101101010",
   "1111100011100101",
   "1111000001000011",
   "1100101000111111",
   "0011000100101111",
   "1100110101110101",
   "1101101010000000",
   "0000010000010110",
   "0011011000011001",
   "0000110011000100",
   "0010010010011011",
   "1100110110010101",
   "0000110001011001",
   "1101111001000011",
   "1111101111000111",
   "0000110001011100",
   "1111010100011000",
   "1101101101101111",
   "0011000010011001",
   "0011010110101101",
   "0010100110110101",
   "1110000101111000",
   "0011101010101011",
   "1101000100111000",
   "1101111101111110",
   "0001001101011000",
   "0000111101011011",
   "1100111101010010",
   "0011010010111110",
   "1101101011100100",
   "1101000001100111",
   "1100110101100000",
   "1110011111101000",
   "1110001000110101",
   "1101110010001101",
   "1111001101010001",
   "1101010011011011",
   "1110101101110110",
   "0010101111001111",
   "0010100001110110",
   "0000001000000001",
   "1101100101000100",
   "0001101010001100",
   "0000001001000111",
   "1111010100100010",
   "1111001000011100",
   "1110101100110111",
   "0010110101000111",
   "0010110000010101");



constant lut_gs_23 : vector_of_std_logic_vector16(0 to 63) := 
  ("1111100111011100",
   "1110100011011111",
   "0010110010111011",
   "1110000001111110",
   "0001110101100111",
   "1111000110000110",
   "1101111010011000",
   "1101110100100110",
   "0011010001110010",
   "0010001101100001",
   "1111010001010000",
   "0001100101111100",
   "0001101011100101",
   "0001100000100000",
   "1101001000010001",
   "0010010100100010",
   "1110110100011111",
   "1110100010000010",
   "1100110111111011",
   "0010111001001011",
   "1100111101001000",
   "1101111000101101",
   "1111100000001010",
   "0011001000010101",
   "0001011111110111",
   "0010010001100100",
   "1101000110110101",
   "0001011101111111",
   "1110000101101111",
   "0000100111001101",
   "0001001100111011",
   "1110101001101000",
   "1101101010001100",
   "0010111101001011",
   "0011001010001100",
   "0010101000110101",
   "1110001010111101",
   "0011010111001111",
   "1101001100001111",
   "1110000101101111",
   "0001111010011111",
   "0001101001100100",
   "1101000100111011",
   "0010111110101000",
   "1101110000010101",
   "1101010100011001",
   "1100111111001110",
   "1110100001101010",
   "1110000100111001",
   "1101110000100010",
   "1110011110000010",
   "1101001111100101",
   "1110100111000111",
   "0010110111101111",
   "0010001101100001",
   "0000110100010000",
   "1101111000101101",
   "0001101111011010",
   "0001000011111011",
   "1110100111011100",
   "1110010010010001",
   "1101111101111011",
   "0010100110001010",
   "0010100001111011");



constant lut_gs_24 : vector_of_std_logic_vector16(0 to 63) := 
  ("1111101010001010",
   "1101111000010111",
   "0010011000100010",
   "1101110100111001",
   "0001111111001110",
   "1110100100110100",
   "1101101100110000",
   "1110000101010111",
   "0010111101001011",
   "0001111110010111",
   "1110100001010011",
   "0001101010110110",
   "0010001001000000",
   "0001101001100111",
   "1101010001010000",
   "0010100001000000",
   "1110001110000010",
   "1110001011111011",
   "1101010010111000",
   "0010100011100101",
   "1101010000100101",
   "1110000101010011",
   "1110101111000011",
   "0010101100011101",
   "0010000000111100",
   "0010001101111100",
   "1101100000101000",
   "0010000001101110",
   "1110001110101010",
   "0001011101111100",
   "0001100100101100",
   "1110000110011010",
   "1101101100101100",
   "0010101011110010",
   "0010110000110111",
   "0010100001000000",
   "1110001100010111",
   "0010110110000001",
   "1101011101100101",
   "1110001010011110",
   "0010010110110000",
   "0010001000100111",
   "1101010111111101",
   "0010100000100111",
   "1101110110100011",
   "1101101101000101",
   "1101010100010011",
   "1110011101010011",
   "1110000000100101",
   "1101110001100110",
   "1101111011010101",
   "1101010110111000",
   "1110011010010101",
   "0010110010111100",
   "0001111010001011",
   "0001011110111010",
   "1110001001100000",
   "0001110111010111",
   "0001110111011111",
   "1110000100101011",
   "1101101011111001",
   "1101100001000111",
   "0010010001101100",
   "0010010000100001");



constant lut_gs_25 : vector_of_std_logic_vector16(0 to 63) := 
  ("1111101111100010",
   "1101011101100001",
   "0001111011000110",
   "1101111001100010",
   "0010001001110110",
   "1110000111100100",
   "1101110010100010",
   "1110010100011100",
   "0010010111101100",
   "0001110100010000",
   "1101110100101000",
   "0001110010100100",
   "0010010110110000",
   "0001110101001110",
   "1101100110000011",
   "0010010111001001",
   "1101110010100010",
   "1101111110011101",
   "1101111010101011",
   "0010000010101011",
   "1101110001111110",
   "1110001111101101",
   "1101111110010011",
   "0010000100010111",
   "0010010000001000",
   "0010000101100000",
   "1110000100010101",
   "0010010111101100",
   "1110010100000011",
   "0010001100010101",
   "0001110110010111",
   "1101101010111110",
   "1101110100101000",
   "0010010000010011",
   "0010001110000010",
   "0010001011111100",
   "1110000111000001",
   "0010001011011000",
   "1101110110101110",
   "1110001000101101",
   "0010011100000100",
   "0010011000110101",
   "1101110100000100",
   "0001111001000001",
   "1101111111011011",
   "1110000111100100",
   "1101110110010101",
   "1110010000000110",
   "1101111110110110",
   "1101110111110110",
   "1101100111001011",
   "1101101000101101",
   "1110001010110010",
   "0010011100100111",
   "0001101000111010",
   "0010000111000001",
   "1110010110101101",
   "0010000011001111",
   "0010100000111101",
   "1101101110001100",
   "1101011100111100",
   "1101011100111100",
   "0001110110110000",
   "0001111100001110");



constant lut_gs_26 : vector_of_std_logic_vector16(0 to 63) := 
  ("1111111011100111",
   "1101011100100000",
   "0001011001111110",
   "1110001000111000",
   "0010001101111100",
   "1101101101000101",
   "1110000100101011",
   "1110011001010111",
   "0001100110000101",
   "0001101010011000",
   "1101010100110001",
   "0010000010110001",
   "0010010000101011",
   "0010001000011001",
   "1110001100101101",
   "0001111110010011",
   "1101100111100110",
   "1101111101011011",
   "1110100110010000",
   "0001011110111010",
   "1110011100111001",
   "1110010000000101",
   "1101010111101111",
   "0001010101010111",
   "0010010010000001",
   "0001111011100000",
   "1110101001001110",
   "0010100001100010",
   "1110001110101010",
   "0010110101010000",
   "0010000100011111",
   "1101011110111100",
   "1110001001011000",
   "0001100101100011",
   "0001011101011110",
   "0001101100100110",
   "1110000001100101",
   "0001010011111011",
   "1110011001001111",
   "1110000010110011",
   "0010001111111010",
   "0010010001110100",
   "1110011010011101",
   "0001010001001010",
   "1110000111011010",
   "1110100100110100",
   "1110011100111001",
   "1101111101101101",
   "1101111001101110",
   "1101111100011000",
   "1101101010010000",
   "1110001011011111",
   "1101110011101100",
   "0001110111101100",
   "0001011110100001",
   "0010100111010011",
   "1110011000001110",
   "0010001111000101",
   "0010110110111000",
   "1101101001000010",
   "1101100001000111",
   "1101101011111001",
   "0001011101000101",
   "0001101101110100");



constant lut_gs_27 : vector_of_std_logic_vector16(0 to 63) := 
  ("0000001010111010",
   "1101101110110100",
   "0000110100011101",
   "1110100111011100",
   "0010010001100100",
   "1101010100011001",
   "1110100111011100",
   "1110011010000100",
   "0000101110110100",
   "0001101000000011",
   "1100111101001000",
   "0010010011000001",
   "0001110101010001",
   "0010011010010100",
   "1110111100000101",
   "0001010011000111",
   "1101110000111110",
   "1110001011100101",
   "1111011000110011",
   "0000110100010000",
   "1111001011110000",
   "1110001101000011",
   "1100110111101011",
   "0000100101010110",
   "0010000000001100",
   "0001110011100001",
   "1111010011010110",
   "0010100010100111",
   "1110000101101111",
   "0011001111101100",
   "0010010001100011",
   "1101011011010010",
   "1110100100001011",
   "0000110101000001",
   "0000101001010100",
   "0001000111010001",
   "1101110110100110",
   "0000011010011010",
   "1111000101100010",
   "1101111100000011",
   "0001101101101111",
   "0001111010101100",
   "1111001010111111",
   "0000100101010110",
   "1110001011001010",
   "1111000110000110",
   "1111001011110000",
   "1101101010111001",
   "1101111000001001",
   "1110000100111001",
   "1101111101101110",
   "1110110110101000",
   "1101011110000101",
   "0001001001011011",
   "0001011110010110",
   "0010111011010010",
   "1110010100101001",
   "0010010110111110",
   "0010111111010101",
   "1101111000010001",
   "1101111101111011",
   "1110010010010001",
   "0000111111000111",
   "0001100000100000");



constant lut_gs_28 : vector_of_std_logic_vector16(0 to 63) := 
  ("0000011011000000",
   "1110010011111101",
   "0000001110101010",
   "1111001111100110",
   "0010010010011011",
   "1101000001100111",
   "1111010100100010",
   "1110010100111100",
   "1111110100110111",
   "0001101010110000",
   "1100110000111001",
   "0010100010111111",
   "0001001010011010",
   "0010101010100101",
   "1111110001111110",
   "0000011101010000",
   "1110001011011111",
   "1110100101110011",
   "0000001011111110",
   "0000001000000001",
   "1111111100111011",
   "1110000101100100",
   "1100100010101011",
   "1111110101101111",
   "0001011111000010",
   "0001101100011111",
   "1111111101110000",
   "0010011010111111",
   "1101111001000011",
   "0011011100110001",
   "0010011011000011",
   "1101100000011001",
   "1111000110001001",
   "0000000000101100",
   "1111110011101110",
   "0000011100100101",
   "1101101010010100",
   "1111100001011100",
   "1111110110000001",
   "1101110011100111",
   "0000111100100000",
   "0001010100000001",
   "1111111111010100",
   "1111111010101011",
   "1110001100100001",
   "1111101000000100",
   "1111111100111011",
   "1101011000011010",
   "1101110111111101",
   "1110001101110001",
   "1110100001010011",
   "1111101000101011",
   "1101001010101111",
   "0000010100000111",
   "0001100101010100",
   "0011000100011011",
   "1110001011010100",
   "0010011100000010",
   "0010111001111011",
   "1110011000000000",
   "1110101100110111",
   "1111001000011100",
   "0000011111110110",
   "0001010111111010");



constant lut_gs_29 : vector_of_std_logic_vector16(0 to 63) := 
  ("0000101000111100",
   "1111000110111111",
   "1111101010010001",
   "1111111100111000",
   "0010010000101110",
   "1100110110101110",
   "0000000110100110",
   "1110001011100111",
   "1110111110000110",
   "0001110001010001",
   "1100110000001000",
   "0010101111101110",
   "0000010101101111",
   "0010110110010100",
   "0000101000101110",
   "1111100011101011",
   "1110110100011000",
   "1111001010000111",
   "0000111011010101",
   "1111011101100010",
   "0000101100001011",
   "1101111011110000",
   "1100011010011001",
   "1111001010000111",
   "0000110010011011",
   "0001100111100100",
   "0000100101100110",
   "0010001101111110",
   "1101101011011101",
   "0011011100101101",
   "0010100000100101",
   "1101101011011101",
   "1111101101011001",
   "1111001101100101",
   "1111000001100011",
   "1111110000001001",
   "1101011111011011",
   "1110101110001000",
   "0000100110011010",
   "1101101011011101",
   "0000000011001000",
   "0000100010011110",
   "0000110010011011",
   "1111010011110101",
   "1110001011100111",
   "0000001001101110",
   "0000101100001011",
   "1101001001101100",
   "1101111001000000",
   "1110010101010100",
   "1111010000101101",
   "0000011100101100",
   "1100111100110111",
   "1111011101100010",
   "0001110001010001",
   "0011000011000010",
   "1101111110111000",
   "0010011101011101",
   "0010101010010010",
   "1111000100101011",
   "1111100111001001",
   "0000000110100110",
   "0000000000000000",
   "0001010100111101");



constant lut_gs_30 : vector_of_std_logic_vector16(0 to 63) := 
  ("0000110001100101",
   "0000000001100001",
   "1111001000110011",
   "0000101010010101",
   "0010001100111111",
   "1100110101100000",
   "0000110111101011",
   "1110000000011011",
   "1110010000011010",
   "0001111001110101",
   "1100111010000001",
   "0010110110001100",
   "1111011110001001",
   "0010111010110011",
   "0001011010000110",
   "1110101110000000",
   "1111100111100001",
   "1111110101101111",
   "0001100010100100",
   "1110111000000101",
   "0001010101010001",
   "1101110010010111",
   "1100011111101100",
   "1110100101110011",
   "1111111111010100",
   "0001100101110100",
   "0001001000001111",
   "0001111111011000",
   "1101100000011001",
   "0011010000101011",
   "0010100001110010",
   "1101111001000011",
   "0000010111011000",
   "1110100000111110",
   "1110010111101100",
   "1111000101111111",
   "1101011000110111",
   "1110000101011010",
   "0001010010000011",
   "1101100101110101",
   "1111001001100101",
   "1111101011111001",
   "0001011111000010",
   "1110110011001001",
   "1110001000110101",
   "0000101010001110",
   "0001010101010001",
   "1101000010001110",
   "1101111010111100",
   "1110011001110111",
   "0000000110011101",
   "0001001101000111",
   "1100110111100010",
   "1110101011111111",
   "0001111111010001",
   "0010111000010101",
   "1101110010101011",
   "0010011010101111",
   "0010010101001100",
   "1111111001011110",
   "0000100100100001",
   "0001000011110001",
   "1111100000001010",
   "0001010111111010");



constant lut_gs_31 : vector_of_std_logic_vector16(0 to 63) := 
  ("0000110010001011",
   "0000111100101000",
   "1110101011011111",
   "0001010011000100",
   "0010000111110111",
   "1100111111001110",
   "0001100001111110",
   "1101110101111111",
   "1101110000111110",
   "0010000010011011",
   "1101001101000101",
   "0010110011110001",
   "1110101010110010",
   "0010110101110111",
   "0010000000001100",
   "1110000011011011",
   "0000011111111010",
   "0000100101010110",
   "0001111110000010",
   "1110011010011111",
   "0001110100011011",
   "1101101100010011",
   "1100110010011110",
   "1110001011100101",
   "1111001010111111",
   "0001101000000011",
   "0001100011011010",
   "0001110010111101",
   "1101011011010010",
   "0010111010100001",
   "0010011110100101",
   "1110000101101111",
   "0001000001010001",
   "1101111111110100",
   "1101111010011000",
   "1110100010000010",
   "1101011001010010",
   "1101101011011110",
   "0001110100011110",
   "1101100100111111",
   "1110010111110001",
   "1110110110100101",
   "0010000000001100",
   "1110011010011111",
   "1110000100111001",
   "0001001000110100",
   "0001110100011011",
   "1101000100111011",
   "1101111101010110",
   "1110011010000100",
   "0000111100101000",
   "0001110100011110",
   "1100111101010101",
   "1110000101010100",
   "0010001100001000",
   "0010100110000111",
   "1101101010001100",
   "0010010011101010",
   "0001111111101101",
   "0000110000111010",
   "0001011100100001",
   "0001110111001001",
   "1111000000111001",
   "0001100000100000");



constant lut_gs_32 : vector_of_std_logic_vector16(0 to 63) := 
  ("0000101000110101",
   "0001110001110111",
   "1110010011001100",
   "0001110010101110",
   "0010000010000101",
   "1101010100010011",
   "0010000000011110",
   "1101101110101000",
   "1101100011011010",
   "0010001001010000",
   "1101100111011110",
   "0010100110101000",
   "1110000010001011",
   "0010100110001010",
   "0010010110001110",
   "1101101001101101",
   "0001011000010101",
   "0001010101010111",
   "0010001011000111",
   "1110000110111110",
   "0010000110110010",
   "1101101100001110",
   "1101010001101001",
   "1101111101011011",
   "1110011010011101",
   "0001101110100100",
   "0001110101010011",
   "0001101011101110",
   "1101011110111100",
   "0010011100011110",
   "0010010111001101",
   "1110001110101010",
   "0001101000001100",
   "1101101101111111",
   "1101101100110000",
   "1110000111101111",
   "1101100010101111",
   "1101100011001101",
   "0010001001111101",
   "1101101010110011",
   "1101110100011111",
   "1110001000010100",
   "0010010010000001",
   "1110001011001011",
   "1110000000100101",
   "0001100100110000",
   "0010000110110010",
   "1101010011110000",
   "1101111111110100",
   "1110010101001010",
   "0001101101101011",
   "0010001110001010",
   "1101001111110101",
   "1101101110001100",
   "0010010101000110",
   "0010001110100001",
   "1101101000100000",
   "0010001000001101",
   "0001101110011000",
   "0001100101100111",
   "0010000111101001",
   "0010011001010001",
   "1110100010111011",
   "0001101101110100");



constant lut_gs_33 : vector_of_std_logic_vector16(0 to 63) := 
  ("0000010111001101",
   "0010011110010011",
   "1101111110010011",
   "0010000011110100",
   "0001111010001001",
   "1101110001111110",
   "0010001101011110",
   "1101101110001100",
   "1101101011100010",
   "0010001111001010",
   "1110000100111010",
   "0010001011111101",
   "1101100111001011",
   "0010001101101001",
   "0010011011011111",
   "1101100110100110",
   "0010001001101011",
   "0010000000000001",
   "0010001010110100",
   "1101111100110001",
   "0010001000100011",
   "1101110110010101",
   "1101111101010101",
   "1101111010000111",
   "1101101111101101",
   "0001110110111010",
   "0001111110111001",
   "0001101001010011",
   "1101101010111110",
   "0001111011000110",
   "0010001010001111",
   "1110010100000011",
   "0010000111011010",
   "1101101111111000",
   "1101101110001100",
   "1101110111011101",
   "1101111000011010",
   "1101101111111000",
   "0010001101110111",
   "1101110110010101",
   "1101100010010000",
   "1101100111101111",
   "0010010100011110",
   "1110000011110001",
   "1101111010100000",
   "0001111011000110",
   "0010001100111001",
   "1101110001011001",
   "1110000100001011",
   "1110001101011100",
   "0010010111010011",
   "0010011001001110",
   "1101101101000011",
   "1101101011100010",
   "0010010110001010",
   "0001110001011100",
   "1101101101101000",
   "0001110110010111",
   "0001100110101001",
   "0010010101000010",
   "0010100010011111",
   "0010100111011010",
   "1110001001010000",
   "0010000000100101");



constant lut_gs_34 : vector_of_std_logic_vector16(0 to 63) := 
  ("1111111001101001",
   "0010111000000110",
   "1101110011100110",
   "0010000110111011",
   "0001110111010011",
   "1110011001001011",
   "0010001001111001",
   "1101101110101000",
   "1110000101111010",
   "0010010000111010",
   "1110100110000010",
   "0001101011001011",
   "1101100011011010",
   "0001100110110001",
   "0010001100110011",
   "1101111000001110",
   "0010110110011111",
   "0010101000101111",
   "0001111010110111",
   "1110000011000010",
   "0001111100001101",
   "1110000100111110",
   "1110101011111000",
   "1110001000001101",
   "1101010100001110",
   "0010000010110001",
   "0001111100111110",
   "0001110010100100",
   "1110000110011010",
   "0001010110000010",
   "0001111011100100",
   "1110001110101010",
   "0010100011101001",
   "1101111111000100",
   "1110000000111101",
   "1101110101010010",
   "1110010011011010",
   "1110001001110110",
   "0010000110000001",
   "1110001010100110",
   "1101101001101101",
   "1101010000110011",
   "0010000100101011",
   "1110001011001011",
   "1101110110000000",
   "0010001101110000",
   "0001111111111100",
   "1110010110000100",
   "1110000111011110",
   "1101111101001111",
   "0010101111111110",
   "0010010001111000",
   "1110010110010001",
   "1101111011001000",
   "0010010001011000",
   "0001010011010001",
   "1110000001010000",
   "0001100000111101",
   "0001100111010100",
   "0010110101000011",
   "0010100011100000",
   "0010011001010001",
   "1101101110010100",
   "0010010100001111");



constant lut_gs_35 : vector_of_std_logic_vector16(0 to 63) := 
  ("1111010100110011",
   "0011000100110010",
   "1101101100010110",
   "0001111110000010",
   "0001110011100001",
   "1111001001101001",
   "0001111000100101",
   "1101110101111111",
   "1110101100111001",
   "0010001100001000",
   "1111001011100011",
   "0000111111111101",
   "1101110000111110",
   "0000111010011110",
   "0001101001100100",
   "1110011001111000",
   "0011010101001000",
   "0011000110001110",
   "0001011010101010",
   "1110010010111001",
   "0001100101100100",
   "1110011110101011",
   "1111100000000110",
   "1110011111111100",
   "1101000010110101",
   "0010010011000001",
   "0001101101000111",
   "0001111111101101",
   "1110101001101000",
   "0000101100110111",
   "0001101111011010",
   "1110000101101111",
   "0010110101000100",
   "1110100000001001",
   "1110100101010110",
   "1110000011111111",
   "1110111000101111",
   "1110110100011111",
   "0001101100111000",
   "1110101001101000",
   "1110000011011011",
   "1101001010011000",
   "0001100001111110",
   "1110011010011111",
   "1101110110000010",
   "0010011110100100",
   "0001100111101011",
   "1111000101011111",
   "1110000111000011",
   "1101101100111111",
   "0010111101001011",
   "0001110110100101",
   "1111001010111111",
   "1110011000100010",
   "0010001010000001",
   "0000110111110011",
   "1110011100100101",
   "0001001010110100",
   "0001101101011101",
   "0011001010001100",
   "0010010001001100",
   "0001110111001001",
   "1101011001110110",
   "0010100100000001");



constant lut_gs_36 : vector_of_std_logic_vector16(0 to 63) := 
  ("1110101100110011",
   "0011000011001110",
   "1101101010001101",
   "0001100111100000",
   "0001110001011010",
   "1111111101001111",
   "0001011001010001",
   "1110000000011011",
   "1111011101110101",
   "0010000100001100",
   "1111110001010110",
   "0000010000000100",
   "1110010000011010",
   "0000001001111111",
   "0000111000100000",
   "1111001001010000",
   "0011100110000100",
   "0011011000101110",
   "0000110000000101",
   "1110101101011001",
   "0001000100101101",
   "1111000000000101",
   "0000010011100100",
   "1111000001011000",
   "1100111101100111",
   "0010100010111111",
   "0001010010100111",
   "0010010000010000",
   "1111010100011000",
   "0000000011111110",
   "0001100101010000",
   "1101111001000011",
   "0010111101100001",
   "1111001100111100",
   "1111010100110110",
   "1110100000000011",
   "1111100011011011",
   "1111101000100000",
   "0001000111010111",
   "1111001111011100",
   "1110101110000000",
   "1101010000011100",
   "0000110010101111",
   "1110110011001001",
   "1101111000010001",
   "0010101010011011",
   "0001000100011001",
   "1111111001001111",
   "1110000101010011",
   "1101011101000001",
   "0010111101011110",
   "0001001100110011",
   "0000000100001111",
   "1111000010010000",
   "0001111111100101",
   "0000011101001100",
   "1111000000011001",
   "0000110001110001",
   "0001111001010011",
   "0011010001110001",
   "0001101100000011",
   "0001000011110001",
   "1101001010111001",
   "0010110000000000");



constant lut_gs_37 : vector_of_std_logic_vector16(0 to 63) := 
  ("1110000110110010",
   "0010110110010100",
   "1101101100010001",
   "0001000101000010",
   "0001110001010001",
   "0000101111010011",
   "0000101111010011",
   "1110001011100111",
   "0000010010100111",
   "0001111010111111",
   "0000010101101111",
   "1111011111110110",
   "1110111110000110",
   "1111011001100110",
   "0000000000000000",
   "0000000000000000",
   "0011101000101111",
   "0011011111000001",
   "0000000000000000",
   "1111010000101101",
   "0000011100101100",
   "1111100111001001",
   "0001000001111010",
   "1111101001100100",
   "1101000011000111",
   "0010101111101110",
   "0000101111010011",
   "0010100000100101",
   "0000000011001000",
   "1111011101011011",
   "0001011110101010",
   "1101101011011101",
   "0010111101010001",
   "0000000000000000",
   "0000001001101110",
   "1111000110111111",
   "0000001111110111",
   "0000011111011101",
   "0000011001100100",
   "1111111001011010",
   "1111100011101011",
   "1101011111011011",
   "1111111100111000",
   "1111010011110101",
   "1101111100001000",
   "0010110000011011",
   "0000011001100100",
   "0000101100001011",
   "1110000010101101",
   "1101010000010010",
   "0010110011001100",
   "0000011001100100",
   "0000111100001001",
   "1111110011001010",
   "0001110100011001",
   "0000000011001000",
   "1111101010010001",
   "0000010101101111",
   "0010000111101110",
   "0011001100110000",
   "0000111001000001",
   "0000000110100110",
   "1101000010101111",
   "0010110110010100");



constant lut_gs_38 : vector_of_std_logic_vector16(0 to 63) := 
  ("1101101000001101",
   "0010100010001010",
   "1101110001010100",
   "0000011001010100",
   "0001110011001010",
   "0001011011000001",
   "1111111110111111",
   "1110010100111100",
   "0001000100101010",
   "0001110010101010",
   "0000110111001101",
   "1110110100000010",
   "1111110100110111",
   "1110101101111101",
   "1111000111100000",
   "0000110110110000",
   "0011011101101010",
   "0011011000101110",
   "1111001111111011",
   "1111111010010110",
   "1111110001000101",
   "0000010001010100",
   "0001100111001011",
   "0000010100111111",
   "1101010000110100",
   "0010110110001100",
   "0000000101101010",
   "0010101100100101",
   "0000110001101101",
   "1110111011001001",
   "0001011100110110",
   "1101100000011001",
   "0010110101000111",
   "0000110011000100",
   "0000111101011011",
   "1111110101011011",
   "0000111010000001",
   "0001010010010100",
   "1111101000010111",
   "0000100100010111",
   "0000011101010000",
   "1101110010101110",
   "1111000111001100",
   "1111111010101011",
   "1110000000101100",
   "0010101111110111",
   "1111101011010101",
   "0001011000111101",
   "1101111111110111",
   "1101001001110100",
   "0010100001110110",
   "1111100010111011",
   "0001101100011000",
   "0000100101011001",
   "0001101011000100",
   "1111101000111000",
   "0000010111000100",
   "1111110110110010",
   "0010010100111011",
   "0010111101010000",
   "1111111110011111",
   "1111001000011100",
   "1101000010011111",
   "0010110101011000");



constant lut_gs_39 : vector_of_std_logic_vector16(0 to 63) := 
  ("1101010110000100",
   "0010001011011010",
   "1101110111111100",
   "1111100111101101",
   "0001110110111101",
   "0001111100000001",
   "1111001101000101",
   "1110011010000100",
   "0001101101101011",
   "0001101101010000",
   "0001010100100001",
   "1110010001000010",
   "0000101110110100",
   "1110001011100010",
   "1110010110011100",
   "0001100110001000",
   "0011000110001110",
   "0011000110001110",
   "1110100101010110",
   "0000100111011101",
   "1111000101100010",
   "0000111011110001",
   "0010000000001000",
   "0000111111111101",
   "1101100011100101",
   "0010110011110001",
   "1111011000100011",
   "0010110000011011",
   "0001011011111000",
   "1110011110101011",
   "0001100000100000",
   "1101011011010010",
   "0010100110001010",
   "0001011111110111",
   "0001101001100100",
   "0000100111011101",
   "0001011101111110",
   "0001111010011111",
   "1110111000101111",
   "0001001100111110",
   "0001010011000111",
   "1110000101100000",
   "1110011000100010",
   "0000100101010110",
   "1110000100111100",
   "0010101000010001",
   "1110111101111100",
   "0001111010101100",
   "1101111101010110",
   "1101001100001111",
   "0010001101100001",
   "1110101111000010",
   "0010001111000110",
   "0001010011000100",
   "0001100101111100",
   "1111001101101101",
   "0001000011010111",
   "1111010101001111",
   "0010011101000111",
   "0010100110000111",
   "1111000011011000",
   "1110010010010001",
   "1101001010111100",
   "0010101100001011");



constant lut_gs_40 : vector_of_std_logic_vector16(0 to 63) := 
  ("1101010100000100",
   "0001110110011100",
   "1101111110101011",
   "1110110100000000",
   "0001111100010100",
   "0010001110111010",
   "1110011110001100",
   "1110011001010111",
   "0010001000100011",
   "0001101100010001",
   "0001101100110100",
   "1101111010011101",
   "0001100110000101",
   "1101110110000011",
   "1101110011001101",
   "0010000111110010",
   "0010100100100010",
   "0010101000101111",
   "1110000101001001",
   "0001010100111001",
   "1110011101011011",
   "0001100011110010",
   "0010001010101010",
   "0001100110111110",
   "1101111000000101",
   "0010100110101000",
   "1110101011000111",
   "0010101001001000",
   "0001111110000000",
   "1110001001001011",
   "0001101001100111",
   "1101011110111100",
   "0010010001101100",
   "0010000000111100",
   "0010001000100111",
   "0001011001000101",
   "0001111000010001",
   "0010010010100100",
   "1110001111001101",
   "0001110000010000",
   "0001111110010011",
   "1110010011100001",
   "1101110110111011",
   "0001010001001010",
   "1110000111111100",
   "0010011001100111",
   "1110010101010011",
   "0010001101101000",
   "1101111011101000",
   "1101011001011000",
   "0001111010001011",
   "1110000011010111",
   "0010011111110001",
   "0001110110111011",
   "0001100110101001",
   "1110110001001001",
   "0001101011111010",
   "1110110001111001",
   "0010011101001000",
   "0010001010010100",
   "1110001110001001",
   "1101101011111001",
   "1101011100010111",
   "0010011010010011");



constant lut_gs_41 : vector_of_std_logic_vector16(0 to 63) := 
  ("1101100001110010",
   "0001100100100011",
   "1110000010000110",
   "1101111111111111",
   "0010000000100101",
   "0010001111100011",
   "1101111000011010",
   "1110010000000110",
   "0010001111101111",
   "0001101110001110",
   "0001111101010111",
   "1101110100110011",
   "0010010011010110",
   "1101110010001001",
   "1101100100100001",
   "0010010101000011",
   "0001111001000001",
   "0010000100010111",
   "1101110000110110",
   "0010000001101101",
   "1101111101101110",
   "0010000100110000",
   "0010000011110100",
   "0010001001010010",
   "1110001001000110",
   "0010010000010011",
   "1110000010101001",
   "0010010111010011",
   "0010010111101100",
   "1101111101010101",
   "0001110101001110",
   "1101101111010100",
   "0001110110110000",
   "0010010000001000",
   "0010010100011110",
   "0010001000101110",
   "0010000100001101",
   "0010011001011010",
   "1101110001011001",
   "0010001110000010",
   "0010011011011111",
   "1110011100000001",
   "1101100100100001",
   "0001111101010111",
   "1110001011001011",
   "0010000110011100",
   "1101110110101110",
   "0010010001110100",
   "1101111101001010",
   "1101101111101101",
   "0001101101010000",
   "1101100110000011",
   "0010011001110011",
   "0010001010110100",
   "0001101111111010",
   "1110010101100101",
   "0010001011110001",
   "1110010000010001",
   "0010010000101100",
   "0001101010011011",
   "1101100001101101",
   "1101011000100110",
   "1101110100001111",
   "0001111101111100");



constant lut_gs_42 : vector_of_std_logic_vector16(0 to 63) := 
  ("1110000011010000",
   "0001011110100001",
   "1110000111111000",
   "1101010010000111",
   "0010000101101111",
   "0010000000011010",
   "1101010111111101",
   "1110000001101001",
   "0010000100110100",
   "0001111001011010",
   "0010001000101011",
   "1101111110001011",
   "0010111001011101",
   "1101111001111111",
   "1101101001110010",
   "0010010010100100",
   "0001001101001110",
   "0001011001000101",
   "1101110001001010",
   "0010100100010101",
   "1101100101101101",
   "0010011111011100",
   "0001101111000000",
   "0010100010001110",
   "1110011010110011",
   "0001101110111001",
   "1101011111011001",
   "0001110100100001",
   "0010100101010000",
   "1101110100010111",
   "0010001000011001",
   "1110001010001000",
   "0001011101000101",
   "0010010010000001",
   "0010001110000101",
   "0010101100011101",
   "0010000110111111",
   "0010001011100001",
   "1101011010100111",
   "0010100010010010",
   "0010100100101110",
   "1110011011001100",
   "1101100110000100",
   "0010100100010101",
   "1110001011101011",
   "0001101000111100",
   "1101100001100000",
   "0010000000011110",
   "1101111111010110",
   "1110010001000111",
   "0001100010001111",
   "1101010110011010",
   "0010000011111010",
   "0010001111000011",
   "0001111110010111",
   "1101111001011010",
   "0010100011101001",
   "1101101011101010",
   "0001111001110011",
   "0001001011001001",
   "1101000111111010",
   "1101011101011001",
   "1110010100000110",
   "0001011110110110");



constant lut_gs_43 : vector_of_std_logic_vector16(0 to 63) := 
  ("1110110011011100",
   "0001011110010110",
   "1110001001000011",
   "1100110000011000",
   "0010001101100100",
   "0001100101100100",
   "1101000100111011",
   "1101110010011111",
   "0001101011100101",
   "0010000101111110",
   "0010010001100011",
   "1110010011001000",
   "0011001111101100",
   "1110010011001000",
   "1101111111110100",
   "0001111010011111",
   "0000011101110000",
   "0000100111011101",
   "1101111111111000",
   "0011000000101110",
   "1101010011110101",
   "0010110101000100",
   "0001010000111101",
   "0010101110010001",
   "1110100101000000",
   "0001000010000100",
   "1101000001011000",
   "0001001001011000",
   "0010100100101110",
   "1101110011111001",
   "0010011010010100",
   "1110101011101110",
   "0000111111000111",
   "0010000000001100",
   "0001111000100101",
   "0011001000010101",
   "0001111001111011",
   "0001101000001111",
   "1101010001101011",
   "0010101010001010",
   "0010010110101001",
   "1110001111001101",
   "1101111101101110",
   "0011000000101110",
   "1110000111000011",
   "0001001000110100",
   "1101010011110101",
   "0001100001111110",
   "1101111111011100",
   "1110111101111100",
   "0001100000011100",
   "1101010001101011",
   "0001011010011011",
   "0010000101101000",
   "0010001101100001",
   "1101011100000000",
   "0010110101000100",
   "1101001101000101",
   "0001011011111000",
   "0000110000001101",
   "1100111011001110",
   "1101111011110101",
   "1110111100101001",
   "0000111000010111");



constant lut_gs_44 : vector_of_std_logic_vector16(0 to 63) := 
  ("1111101100111111",
   "0001100101010100",
   "1110000111111010",
   "1100011011000101",
   "0010010100110001",
   "0000111111110001",
   "1100111101010010",
   "1101100011000110",
   "0001000100111110",
   "0010010011111100",
   "0010010110000111",
   "1110110011101101",
   "0011010111110110",
   "1110111000101001",
   "1110100101111010",
   "0001010010010100",
   "1111101111111111",
   "1111110101011011",
   "1110011101110000",
   "0011010010101001",
   "1101001010101000",
   "0011000010011101",
   "0000101010101001",
   "0010110000001000",
   "1110101001001111",
   "0000001111101111",
   "1100101101000010",
   "0000010111010101",
   "0010011010101011",
   "1101111000000111",
   "0010101010100101",
   "1111010100000011",
   "0000011111110110",
   "0001011111000010",
   "0001010100010110",
   "0011011000011001",
   "0001100000010001",
   "0000110110011011",
   "1101010011000110",
   "0010101000111001",
   "0001110101010110",
   "1101111101000110",
   "1110100110001110",
   "0011010010101001",
   "1110000000010111",
   "0000100101010010",
   "1101001111100100",
   "0000110111101011",
   "1101111111100011",
   "1111110000010001",
   "0001100101000000",
   "1101011000000010",
   "0000100100110110",
   "0001101101010000",
   "0010011100111010",
   "1101000010011011",
   "0010111101100001",
   "1100110101000101",
   "0000110110101001",
   "0000010111011100",
   "1100111100110010",
   "1110101101001100",
   "1111101000111100",
   "0000001111001111");



constant lut_gs_45 : vector_of_std_logic_vector16(0 to 63) := 
  ("0000101000111100",
   "0001110001010001",
   "1110000101000001",
   "1100010011110100",
   "0010011001111111",
   "0000010010111111",
   "1100111111111111",
   "1101010110100010",
   "0000010101101111",
   "0010100000100101",
   "0010010110110111",
   "1111011100101110",
   "0011010011000000",
   "1111100110011100",
   "1111010111010010",
   "0000011111011101",
   "1111000110111111",
   "1111000110111111",
   "1111000111110011",
   "0011011000110001",
   "1101001001101100",
   "0011000110111110",
   "0000000000000000",
   "0010101001011110",
   "1110100111100110",
   "1111011100101110",
   "1100100100000111",
   "1111100011010100",
   "0010001010110110",
   "1101111110111000",
   "0010110110010100",
   "0000000000000000",
   "0000000000000000",
   "0000110010011011",
   "0000100101100110",
   "0011011011111001",
   "0000111100001001",
   "1111111100111000",
   "1101011100010011",
   "0010100000100101",
   "0001000101000010",
   "1101101001001001",
   "1111011010011010",
   "0011011000110001",
   "1101111001000000",
   "0000000000000000",
   "1101010011011010",
   "0000000110100110",
   "1101111111100101",
   "0000100011010010",
   "0001101110001001",
   "1101100110000001",
   "1111101010010001",
   "0001001000001010",
   "0010101001011110",
   "1100110000001000",
   "0010111101010001",
   "1100100110011011",
   "0000001100110110",
   "0000000000000000",
   "1101001001101100",
   "1111101010010001",
   "0000010101101111",
   "1111100110011100");



constant lut_gs_46 : vector_of_std_logic_vector16(0 to 63) := 
  ("0001011111100110",
   "0001111111010001",
   "1110000001010000",
   "1100011011000101",
   "0010011011111000",
   "1111100011101111",
   "1101001011000100",
   "1101001111111000",
   "1111100011100101",
   "0010101000111001",
   "0010010100011100",
   "0000001010010011",
   "0011000011010101",
   "0000010111101001",
   "0000001110000010",
   "1111101000100000",
   "1110100101011111",
   "1110100000000011",
   "1111111001110010",
   "0011010010101001",
   "1101010000000000",
   "0011000010011101",
   "1111010101010111",
   "0010011100111010",
   "1110100000110100",
   "1110101110010001",
   "1100100111100111",
   "1110110010111001",
   "0001111001100111",
   "1110000101111000",
   "0010111010110011",
   "0000101011111101",
   "1111100000001010",
   "1111111111010100",
   "1111110001101001",
   "0011010010111110",
   "0000010000010110",
   "1111000011100000",
   "1101101010000000",
   "0010010011111100",
   "0000001011011110",
   "1101011000010110",
   "0000010011110011",
   "0011010010101001",
   "1101110010100001",
   "1111011010101110",
   "1101011101010110",
   "1111010100100010",
   "1101111111100011",
   "0001010001101111",
   "0001111001100000",
   "1101110111010110",
   "1110110010101000",
   "0000011001101000",
   "0010110000001000",
   "1100101000011111",
   "0010110101000111",
   "1100100011100011",
   "1111100001101110",
   "1111101000100100",
   "1101011101110110",
   "0000101010010001",
   "0000111111100111",
   "1111000001000011");



constant lut_gs_47 : vector_of_std_logic_vector16(0 to 63) := 
  ("0010001001101001",
   "0010001100001000",
   "1101111101100101",
   "1100110000011000",
   "0010011001001010",
   "1110110110101000",
   "1101011011111111",
   "1101010001101111",
   "1110110100011111",
   "0010101010001010",
   "0010001111101011",
   "0000111000010111",
   "0010101011100111",
   "0001000111010001",
   "0001000011111011",
   "1110110100011111",
   "1110001101101100",
   "1110000011111111",
   "0000101110110100",
   "0011000000101110",
   "1101011011111111",
   "0010110101000100",
   "1110101111000011",
   "0010001101100001",
   "1110010110000110",
   "1110001001011011",
   "1100110111101011",
   "1110001011100010",
   "0001101011010111",
   "1110001010111101",
   "0010110101110111",
   "0001010100010010",
   "1111000000111001",
   "1111001010111111",
   "1110111110001011",
   "0010111110101000",
   "1111100000001010",
   "1110010010010001",
   "1101111000101101",
   "0010000101111110",
   "1111001111000110",
   "1101001111100101",
   "0001001011100010",
   "0011000000101110",
   "1101101110011100",
   "1110110111001100",
   "1101101010111001",
   "1110100111011100",
   "1101111111011100",
   "0001110110100101",
   "0010000100100001",
   "1110000111100111",
   "1110000101100001",
   "1111100101100110",
   "0010101110010001",
   "1100101110001110",
   "0010100110001010",
   "1100101110001110",
   "1110111000100010",
   "1111001111110011",
   "1101110100100110",
   "0001100100001000",
   "0001100011011011",
   "1110100010000010");



constant lut_gs_48 : vector_of_std_logic_vector16(0 to 63) := 
  ("0010100001001100",
   "0010010101000110",
   "1101111010111101",
   "1101010010000111",
   "0010010000110100",
   "1110001111101011",
   "1101101111111101",
   "1101011101110010",
   "1110001110000010",
   "0010100010010010",
   "0010001001011101",
   "0001100011000011",
   "0010001110101110",
   "0001110000110011",
   "0001110011010011",
   "1110001001110110",
   "1110000001001001",
   "1101110101010010",
   "0001100001111000",
   "0010100100010101",
   "1101101011110001",
   "0010011111011100",
   "1110010001000000",
   "0001111110010111",
   "1110001000110110",
   "1101110010010100",
   "1101010011100011",
   "1101110001110110",
   "0001100011100110",
   "1110001100010111",
   "0010100110001010",
   "0001110101111000",
   "1110100010111011",
   "1110011010011101",
   "1110010000011100",
   "0010100000100111",
   "1110101111000011",
   "1101110000000110",
   "1110000101010011",
   "0001111001011010",
   "1110010110001101",
   "1101010010101100",
   "0001111011011011",
   "0010100100010101",
   "1101101101111000",
   "1110010111000100",
   "1101111001100001",
   "1110000100101011",
   "1101111111010110",
   "0010001101101100",
   "0010001100111110",
   "1110010011000011",
   "1101101001010000",
   "1110110000010010",
   "0010100010001110",
   "1101000010110101",
   "0010010001101100",
   "1101000111000001",
   "1110010100001010",
   "1110110100110111",
   "1110001001100100",
   "0010001111110001",
   "0001111110110000",
   "1110001011111011");



constant lut_gs_49 : vector_of_std_logic_vector16(0 to 63) := 
  ("0010100100111101",
   "0010010110001010",
   "1101111100001101",
   "1101111011101001",
   "0010000100010111",
   "1101110100000100",
   "1110000110011100",
   "1101110010010111",
   "1101110010100010",
   "0010010010011000",
   "0010000000100101",
   "0010000100111100",
   "0001101101000101",
   "0010010010111101",
   "0010010101100111",
   "1101101111111000",
   "1110000010110011",
   "1101110111011101",
   "0010001100010101",
   "0010000001101101",
   "1101111111011011",
   "0010000100110000",
   "1101111100001100",
   "0001101111111010",
   "1101111000011011",
   "1101101101110011",
   "1101110111010010",
   "1101101011001001",
   "0001100010010010",
   "1110000111000001",
   "0010001101101001",
   "0010010000101100",
   "1110000100111010",
   "1101101111101101",
   "1101101010011001",
   "0001111101010111",
   "1101111110010011",
   "1101100011111100",
   "1110001111101101",
   "0001101110001110",
   "1101100011111110",
   "1101100110000011",
   "0010011100100111",
   "0010000001101101",
   "1101110011100000",
   "1101111101111010",
   "1110001001000110",
   "1101110010100010",
   "1110000001100000",
   "0010010110100100",
   "0010010011100000",
   "1110011001010111",
   "1101011111100110",
   "1101111011101001",
   "0010001001010010",
   "1101101000010100",
   "0001110110110000",
   "1101101010111110",
   "1101111000111111",
   "1110011001111011",
   "1110011011011101",
   "0010100101001001",
   "0010001110000010",
   "1101111110011101");



constant lut_gs_50 : vector_of_std_logic_vector16(0 to 63) := 
  ("0010001111101111",
   "0010010001011000",
   "1101111010111101",
   "1110110000010010",
   "0001110001000000",
   "1101100010101111",
   "1110011010010101",
   "1110010101010011",
   "1101100111100110",
   "0001110011111110",
   "0001111000100110",
   "0010100010011011",
   "0001001111010101",
   "0010101001001000",
   "0010101011000001",
   "1101100011001101",
   "1110001011111011",
   "1110000111101111",
   "0010110001010101",
   "0001010100111001",
   "1110010010001100",
   "0001100011110010",
   "1101110101010110",
   "0001100110101001",
   "1101101100111111",
   "1101111001111111",
   "1110100110111011",
   "1101110001110110",
   "0001101110011000",
   "1110000001100101",
   "0001100110110001",
   "0010100001000100",
   "1101101010100101",
   "1101010100001110",
   "1101010001010000",
   "0001010100111001",
   "1101010111101111",
   "1101101001010000",
   "1110010000000101",
   "0001101100010001",
   "1101000010110101",
   "1110000111000101",
   "0010101111001101",
   "0001010100111001",
   "1101111100011000",
   "1101101010000111",
   "1110010101001010",
   "1101101100110000",
   "1101111111010110",
   "0010001001110000",
   "0010010000111010",
   "1110010011000011",
   "1101101100010111",
   "1101010010000111",
   "0001100110111110",
   "1110011001111011",
   "0001011101000101",
   "1110011110010101",
   "1101100101101001",
   "1101111001011010",
   "1110100001011111",
   "0010100011111110",
   "0010010011110010",
   "1101111101011011");



constant lut_gs_51 : vector_of_std_logic_vector16(0 to 63) := 
  ("0001100110001011",
   "0010001010000001",
   "1101111101100101",
   "1111100101100110",
   "0001010100100001",
   "1101011001010010",
   "1110100111000111",
   "1110111101111100",
   "1101110000111110",
   "0001001111000101",
   "0001110100110110",
   "0010110011110001",
   "0000110000001101",
   "0010110000011011",
   "0010110101101000",
   "1101101011011110",
   "1110100010000010",
   "1110100010000010",
   "0011001000000101",
   "0000100111011101",
   "1110011111100000",
   "0000111011110001",
   "1101111111111000",
   "0001100101111100",
   "1101100001011011",
   "1110010011001000",
   "1111011000100011",
   "1110001011100010",
   "0001111111101101",
   "1101110110100110",
   "0000111010011110",
   "0010100100101110",
   "1101010111101111",
   "1101000010110101",
   "1101001000010001",
   "0000100111011101",
   "1100110111101011",
   "1110000101100001",
   "1110001101000011",
   "0001101101010000",
   "1100101110001110",
   "1110110001001000",
   "0010110101101000",
   "0000100111011101",
   "1110000100111001",
   "1101011001110110",
   "1110011010000100",
   "1101111010011000",
   "1101111111011100",
   "0001101110111110",
   "0010001100001000",
   "1110000111100111",
   "1110010000001011",
   "1100110000011000",
   "0000111111111101",
   "1111010001001100",
   "0000111111000111",
   "1111010110101100",
   "1101010111111100",
   "1101011100000000",
   "1110100001101010",
   "0010001111000110",
   "0010010011101101",
   "1110001011100101");



constant lut_gs_52 : vector_of_std_logic_vector16(0 to 63) := 
  ("0000101101111001",
   "0001111111100101",
   "1110000001010000",
   "0000011001101000",
   "0000110010010001",
   "1101011000110111",
   "1110101101110110",
   "1111101011010101",
   "1110001011011111",
   "0000100100000011",
   "0001110011011111",
   "0010111011001000",
   "0000010010100000",
   "0010101100100101",
   "0010110100011111",
   "1110000101011010",
   "1111000001000011",
   "1111000101111111",
   "0011010010000101",
   "1111111010010110",
   "1110101000000110",
   "0000010001010100",
   "1110011000110101",
   "0001101011000100",
   "1101011001010010",
   "1110111000101001",
   "0000001010100101",
   "1110110010111001",
   "0010010101001100",
   "1101101010010100",
   "0000001001111111",
   "0010011111100111",
   "1101001011001110",
   "1100111101100111",
   "1101001011110101",
   "1111111010010110",
   "1100100010101011",
   "1110110010101000",
   "1110000101100100",
   "0001110010101010",
   "1100101000011111",
   "1111100010100110",
   "0010101111100100",
   "1111111010010110",
   "1110001101110001",
   "1101001111110101",
   "1110011001110111",
   "1110010111101100",
   "1101111111100011",
   "0001000111000011",
   "0010000100001100",
   "1101110111010110",
   "1111000011110100",
   "1100011011000101",
   "0000010100111111",
   "0000001011001001",
   "0000011111110110",
   "0000010001001110",
   "1101010001110111",
   "1101000010011011",
   "1110011010101100",
   "0001100111011100",
   "0010001101101001",
   "1110100101110011");



constant lut_gs_53 : vector_of_std_logic_vector16(0 to 63) := 
  ("1111101110101110",
   "0001110100011001",
   "1110000101000001",
   "0001001000001010",
   "0000001100000001",
   "1101011111011011",
   "1110101110001011",
   "0000011001100100",
   "1110110100011000",
   "1111110110010010",
   "0001110100011001",
   "0010111001011100",
   "1111110110010010",
   "0010100000100101",
   "0010101010010010",
   "1110101110001000",
   "1111100110011100",
   "1111110000001001",
   "0011001111111000",
   "1111010000101101",
   "1110101011000011",
   "1111100111001001",
   "1110111110000110",
   "0001110100011001",
   "1101010101101110",
   "1111100110011100",
   "0000111001000001",
   "1111100011010100",
   "0010101010010010",
   "1101011111011011",
   "1111011001100110",
   "0010010100100011",
   "1101000101110111",
   "1101000011000111",
   "1101011000110110",
   "1111010000101101",
   "1100011010011001",
   "1111101010010001",
   "1101111011110000",
   "0001111010111111",
   "1100110000001000",
   "0000010110011100",
   "0010100000100101",
   "1111010000101101",
   "1110010101010100",
   "1101001100011101",
   "1110010101010100",
   "1111000001100011",
   "1101111111100101",
   "0000010110011100",
   "0001111010111111",
   "1101100110000001",
   "0000000000000000",
   "1100010011110100",
   "1111101001100100",
   "0001000001111010",
   "0000000000000000",
   "0001001000001010",
   "1101010010100110",
   "1100110000001000",
   "1110001110101111",
   "0000110010011011",
   "0010000100010000",
   "1111001010000111");



constant lut_gs_54 : vector_of_std_logic_vector16(0 to 63) := 
  ("1110110001101011",
   "0001101011000100",
   "1110000111111010",
   "0001101101010000",
   "1111100100000000",
   "1101101010010100",
   "1110101000011010",
   "0001000100011001",
   "1111100111100001",
   "1111001001101100",
   "0001110111001011",
   "0010110000010101",
   "1111011011001110",
   "0010010000010000",
   "0010011010101000",
   "1111100001011100",
   "0000001111001111",
   "0000011100100101",
   "0011000011000001",
   "1110101101011001",
   "1110101000000110",
   "1111000000000101",
   "1111101100011100",
   "0001111111100101",
   "1101010111100111",
   "0000010111101001",
   "0001011111111101",
   "0000010111010101",
   "0010111001111011",
   "1101011000110111",
   "1110101101111101",
   "0010000110111101",
   "1101001000001111",
   "1101010000110100",
   "1101101011001001",
   "1110101101011001",
   "1100011111101100",
   "0000100100110110",
   "1101110010010111",
   "0010000100001100",
   "1101000010011011",
   "0001000111000011",
   "0010001101010010",
   "1110101101011001",
   "1110011001110111",
   "1101001111110101",
   "1110001101110001",
   "1111110011101110",
   "1101111111100011",
   "1111100010100110",
   "0001110010101010",
   "1101011000000010",
   "0000111100001100",
   "1100011011000101",
   "1111000001011000",
   "0001101111100110",
   "1111100000001010",
   "0001110101101010",
   "1101011000111110",
   "1100101000011111",
   "1110000000101111",
   "1111110110111001",
   "0001111010011100",
   "1111110101101111");



constant lut_gs_55 : vector_of_std_logic_vector16(0 to 63) := 
  ("1101111111100110",
   "0001100101111100",
   "1110001001000011",
   "0010000101101000",
   "1110111100101001",
   "1101110110100110",
   "1110011101011010",
   "0001100111101011",
   "0000011111111010",
   "1110100010000001",
   "0001111011000111",
   "0010100001111011",
   "1111000000111001",
   "0001111111101101",
   "0010001001011010",
   "0000011010011010",
   "0000111000010111",
   "0001000111010001",
   "0010101101101101",
   "1110010010111001",
   "1110011111100000",
   "1110011110101011",
   "0000011111111010",
   "0010001010000001",
   "1101011111100011",
   "0001000111010001",
   "0001111100000001",
   "0001001001011000",
   "0010111111010101",
   "1101011001010010",
   "1110001011100010",
   "0001111010010001",
   "1101010010100010",
   "1101100011100101",
   "1101111110001100",
   "1110010010111001",
   "1100110010011110",
   "0001011010011011",
   "1101101100010011",
   "0010001100001000",
   "1101011100000000",
   "0001101110111110",
   "0001111010100000",
   "1110010010111001",
   "1110011010000100",
   "1101011001110110",
   "1110000100111001",
   "0000101001010100",
   "1101111111011100",
   "1110110001001000",
   "0001101101010000",
   "1101010001101011",
   "0001101111110101",
   "1100110000011000",
   "1110011111111100",
   "0010001111000010",
   "1111000000111001",
   "0010010100100010",
   "1101100011100010",
   "1100101110001110",
   "1101110011111000",
   "1110111100000101",
   "0001110010111101",
   "0000100101010110");



constant lut_gs_56 : vector_of_std_logic_vector16(0 to 63) := 
  ("1101011111110111",
   "0001100110101001",
   "1110000111111000",
   "0010001111000011",
   "1110011000010010",
   "1110000001100101",
   "1110001110011110",
   "0001111111111100",
   "0001011000010101",
   "1110000010011110",
   "0001111111011011",
   "0010010000100001",
   "1110100111000111",
   "0001110010100100",
   "0001111010001111",
   "0001010011111011",
   "0001011110110110",
   "0001101100100110",
   "0010010010011101",
   "1110000011000010",
   "1110010010001100",
   "1110000100111110",
   "0001010100001000",
   "0010010001011000",
   "1101101101110001",
   "0001110000110011",
   "0010001010101110",
   "0001110100100001",
   "0010110110111000",
   "1101100010101111",
   "1101110110000011",
   "0001110001010110",
   "1101100100100000",
   "1101111000000101",
   "1110001101111010",
   "1110000011000010",
   "1101010001101001",
   "0010000011111010",
   "1101101100001110",
   "0010010000111010",
   "1101111001011010",
   "0010001001110000",
   "0001101100011111",
   "1110000011000010",
   "1110010101001010",
   "1101101010000111",
   "1101111100011000",
   "0001011101011110",
   "1101111111010110",
   "1110000111000101",
   "0001101100010001",
   "1101010110011010",
   "0010010011101001",
   "1101010010000111",
   "1110001000001101",
   "0010011100100110",
   "1110100010111011",
   "0010100001000000",
   "1101110000101110",
   "1101000010110101",
   "1101101010111010",
   "1110001000100001",
   "0001101111111011",
   "0001010101010111");



constant lut_gs_57 : vector_of_std_logic_vector16(0 to 63) := 
  ("1101010101000110",
   "0001101111111010",
   "1110000010000110",
   "0010000110011110",
   "1101111011010000",
   "1110000111000001",
   "1101111111011011",
   "0010001100111001",
   "0010001001101011",
   "1101101111010100",
   "0010000001001010",
   "0010000000100101",
   "1110001011111010",
   "0001101001010011",
   "0001110001111111",
   "0010000111000001",
   "0001111101111100",
   "0010000111100110",
   "0001110101110010",
   "1101111100110001",
   "1110000011110010",
   "1101110110010101",
   "0010000111000001",
   "0010010110001010",
   "1101111111111111",
   "0010001110100111",
   "0010001000100011",
   "0010010111010011",
   "0010011100100111",
   "1101110100000100",
   "1101110010001001",
   "0001101011111101",
   "1101111111100110",
   "1110001101011100",
   "1110011001010111",
   "1110000001000111",
   "1101111101010101",
   "0010011001110011",
   "1101110110010101",
   "0010010011100000",
   "1110011001111011",
   "0010010010001101",
   "0001101000010101",
   "1110000001000111",
   "1110001001000110",
   "1101111101111010",
   "1101110111110110",
   "0010001110000010",
   "1110000001100000",
   "1101100110000011",
   "0001101110001110",
   "1101101010011001",
   "0010100100110000",
   "1101111011101001",
   "1101111010000111",
   "0010011000110101",
   "1110000100111010",
   "0010010111001001",
   "1101111100110001",
   "1101100011111110",
   "1101100101011111",
   "1101100011011001",
   "0001110000010011",
   "0010000010001100");



constant lut_gs_58 : vector_of_std_logic_vector16(0 to 63) := 
  ("1101100101010111",
   "0001111110010111",
   "1101111110101011",
   "0001110011001100",
   "1101100100100000",
   "1110001100010111",
   "1101101111011111",
   "0010000110110010",
   "0010110110011111",
   "1101100110100111",
   "0010000110010010",
   "0001110001100010",
   "1101110010101110",
   "0001101011101110",
   "0001101011100001",
   "0010110010010010",
   "0010011010010011",
   "0010011101010001",
   "0001010011000100",
   "1110000110111110",
   "1101101111011111",
   "1101101100001110",
   "0010110010000101",
   "0010010101000110",
   "1110011000010110",
   "0010100101011001",
   "0001111000010001",
   "0010101001001000",
   "0001110011110001",
   "1110001111101011",
   "1101111001111111",
   "0001110001010110",
   "1110011100000001",
   "1110011110100001",
   "1110011100011010",
   "1110001010101101",
   "1110101011111000",
   "0010011111110001",
   "1110000100111110",
   "0010001100111110",
   "1110110100110111",
   "0010001001111101",
   "0001101000100011",
   "1110001010101101",
   "1101111001100001",
   "1110010111000100",
   "1101110001100110",
   "0010110000110111",
   "1101111111010110",
   "1101010010101100",
   "0001111001011010",
   "1110000111000101",
   "0010011010011111",
   "1110110000010010",
   "1101111101011011",
   "0001111101110101",
   "1101101010100101",
   "0001111110010011",
   "1110001000110110",
   "1110010110001101",
   "1101101010111010",
   "1101001100110111",
   "0001111010101101",
   "0010101010100110");



constant lut_gs_59 : vector_of_std_logic_vector16(0 to 63) := 
  ("1110001100100001",
   "0010001101100001",
   "1101110111111100",
   "0001010000111101",
   "1101010010100010",
   "1110001010111101",
   "1101011110000101",
   "0001110100011011",
   "0011010101001000",
   "1101100100111111",
   "0010000111110111",
   "0001100010100110",
   "1101011111010101",
   "0001110010111101",
   "0001101101011101",
   "0011010101001000",
   "0010101100001011",
   "0010100110101110",
   "0000110010010011",
   "1110011010011111",
   "1101011110000101",
   "1101101100010011",
   "0011001111101000",
   "0010001100001000",
   "1110111000100010",
   "0010101110010101",
   "0001011101111110",
   "0010110000011011",
   "0001000001110101",
   "1110110110101000",
   "1110010011001000",
   "0001111010010001",
   "1110111110101111",
   "1110100111000111",
   "1110010100101001",
   "1110011100100110",
   "1111100000000110",
   "0010001111000110",
   "1110011110101011",
   "0010000100100001",
   "1111001111110011",
   "0001110100011110",
   "0001110010111010",
   "1110011100100110",
   "1101101010111001",
   "1110110111001100",
   "1101110000100010",
   "0011001010001100",
   "1101111111011100",
   "1101001111100101",
   "0010000101111110",
   "1110110001001000",
   "0001111100100101",
   "1111100101100110",
   "1110001011100101",
   "0001010101001110",
   "1101010111101111",
   "0001010011000111",
   "1110010110000110",
   "1111001111000110",
   "1101110011111000",
   "1101000010110001",
   "0010000111010011",
   "0011000111010001");



constant lut_gs_60 : vector_of_std_logic_vector16(0 to 63) := 
  ("1111000100111101",
   "0010011100111010",
   "1101110001010100",
   "0000100101101110",
   "1101001000001111",
   "1110000101111000",
   "1101001111101011",
   "0001010101010001",
   "0011100110000100",
   "1101101010110001",
   "0010001000000011",
   "0001010111100110",
   "1101010000111110",
   "0001111111011000",
   "0001110100010111",
   "0011101011000000",
   "0010110101011000",
   "0010100111001001",
   "0000010010001100",
   "1110111000000101",
   "1101001111101011",
   "1101110010010111",
   "0011011111111111",
   "0001111111010001",
   "1111011100110010",
   "0010101100111010",
   "0000111010000001",
   "0010101100100101",
   "0000001001011011",
   "1111100011101111",
   "1110111000101001",
   "0010000110111101",
   "1111100011101100",
   "1110101000111010",
   "1110000110011001",
   "1110110111110001",
   "0000010011100100",
   "0001101100011000",
   "1111000000000101",
   "0001111001100000",
   "1111101000100100",
   "0001010010000011",
   "0010000010100110",
   "1110110111110001",
   "1101011101010110",
   "1111011010101110",
   "1101110010001101",
   "0011010110101101",
   "1101111111100011",
   "1101011000010110",
   "0010010011111100",
   "1111100010100110",
   "0001001101000100",
   "0000011001101000",
   "1110100101110011",
   "0000100001110111",
   "1101001011001110",
   "0000011101010000",
   "1110100000110100",
   "0000001011011110",
   "1110000000101111",
   "1101000101110000",
   "0010010110000000",
   "0011011000100100");



constant lut_gs_61 : vector_of_std_logic_vector16(0 to 63) := 
  ("0000000110011011",
   "0010101001011110",
   "1101101100010001",
   "1111110110010010",
   "1101000101110111",
   "1101111110111000",
   "1101000110100100",
   "0000101100001011",
   "0011101000101111",
   "1101110101001010",
   "0010000111000000",
   "0001010001110101",
   "1101001000111111",
   "0010001101111110",
   "0001111110000000",
   "0011110010011100",
   "0010110110010100",
   "0010100000100101",
   "1111110011001010",
   "1111011101100010",
   "1101000110100100",
   "1101111011110000",
   "0011100010011111",
   "0001110001010001",
   "0000000011001000",
   "0010100011101101",
   "0000001111110111",
   "0010100000100101",
   "1111010000101101",
   "0000010010111111",
   "1111100110011100",
   "0010010100100011",
   "0000001000111001",
   "1110100100011110",
   "1101110101001010",
   "1111011010011010",
   "0001000001111010",
   "0000111100001001",
   "1111100111001001",
   "0001101110001001",
   "0000000000000000",
   "0000100110011010",
   "0010010011101111",
   "1111011010011010",
   "1101010011011010",
   "0000000000000000",
   "1101110101111000",
   "0011010110011101",
   "1101111111100101",
   "1101101001001001",
   "0010100000100101",
   "0000010110011100",
   "0000010010100111",
   "0001001000001010",
   "1111001010000111",
   "1111101010010001",
   "1101000101110111",
   "1111100011101011",
   "1110100111100110",
   "0001000101000010",
   "1110001110101111",
   "1101010010100110",
   "0010100011101101",
   "0011011101011101");



constant lut_gs_62 : vector_of_std_logic_vector16(0 to 63) := 
  ("0001000111001110",
   "0010110000001000",
   "1101101010001101",
   "1111001000000000",
   "1101001011001110",
   "1101111000000111",
   "1101000100111000",
   "1111111100111011",
   "0011011101101010",
   "1110000000111101",
   "0010000101000100",
   "0001010010001010",
   "1101001000100100",
   "0010011010111111",
   "0010000111100101",
   "0011101011000000",
   "0010110000000000",
   "0010010101101100",
   "1111010101011110",
   "0000001000000001",
   "1101000100111000",
   "1110000101100100",
   "0011010111100101",
   "0001100101010100",
   "0000101001010011",
   "0010010110000000",
   "1111100011011011",
   "0010010000010000",
   "1110011110010100",
   "0000111111110001",
   "0000010111101001",
   "0010011111100111",
   "0000101100100001",
   "1110011011000100",
   "1101100101010101",
   "0000000010010000",
   "0001100111001011",
   "0000000100001111",
   "0000010001010100",
   "0001100101000000",
   "0000010111011100",
   "1111110110000001",
   "0010100001111001",
   "0000000010010000",
   "1101001111100100",
   "0000100101010010",
   "1101111010100111",
   "0011001010100110",
   "1101111111100011",
   "1101111101000110",
   "0010101000111001",
   "0001000111000011",
   "1111010101011010",
   "0001101101010000",
   "1111110101101111",
   "1110110101100110",
   "1101001000001111",
   "1110101110000000",
   "1110101001001111",
   "0001110101010110",
   "1110011010101100",
   "1101100101000100",
   "0010101100111010",
   "0011010101110110");



constant lut_gs_63 : vector_of_std_logic_vector16(0 to 63) := 
  ("0001111101101100",
   "0010101110010001",
   "1101101100010110",
   "1110100000001001",
   "1101010111101111",
   "1101110011111001",
   "1101001100001111",
   "1111001011110000",
   "0011000110001110",
   "1110001010111101",
   "0010000010101010",
   "0001011000111001",
   "1101010000011011",
   "0010100010100111",
   "0010001110001101",
   "0011010101001000",
   "0010100100000001",
   "0010001001011010",
   "1110111001010011",
   "0000110100010000",
   "1101001100001111",
   "1110001101000011",
   "0011000000101110",
   "0001011110010110",
   "0001001100111110",
   "0010000111010011",
   "1110111000101111",
   "0001111111101101",
   "1101111000100001",
   "0001100101100100",
   "0001000111010001",
   "0010100100101110",
   "0001001100111011",
   "1110001110100000",
   "1101011011010010",
   "0000101100101010",
   "0010000000001000",
   "1111001010111111",
   "0000111011110001",
   "0001100000011100",
   "0000110000001101",
   "1111000101100010",
   "0010101000110101",
   "0000101100101010",
   "1101010011110101",
   "0001001000110100",
   "1101111111011100",
   "0010110101000001",
   "1101111111011100",
   "1110001111001101",
   "0010101010001010",
   "0001101110111110",
   "1110011101111111",
   "0010000101101000",
   "0000100101010110",
   "1110001010101111",
   "1101010010100010",
   "1110000011011011",
   "1110100101000000",
   "0010010110101001",
   "1110100001101010",
   "1101111000101101",
   "0010101110010101",
   "0011000010011011");



constant lut_gs_64 : vector_of_std_logic_vector16(0 to 63) := 
  ("0010100001101000",
   "0010100010001110",
   "1101110011100110",
   "1110000011010000",
   "1101101010100101",
   "1101110100010111",
   "1101011101100101",
   "1110011100111001",
   "0010100100100010",
   "1110010000100011",
   "0010000000001100",
   "0001100101101011",
   "1101100000110001",
   "0010100001100010",
   "0010001111011000",
   "0010110010010010",
   "0010010100001111",
   "0001111110011011",
   "1110011110111111",
   "0001011110111010",
   "1101011101100101",
   "1110010000000101",
   "0010100000001001",
   "0001011110100001",
   "0001101100000011",
   "0001111010101101",
   "1110010011011010",
   "0001110010100100",
   "1101100100001011",
   "0010000000011010",
   "0001110000110011",
   "0010100001000100",
   "0001101000111000",
   "1110000000101110",
   "1101011010110000",
   "0001010110110010",
   "0010001010101010",
   "1110010110010001",
   "0001100011110010",
   "0001100010001111",
   "0001001011001001",
   "1110011001001111",
   "0010100101001100",
   "0001010110110010",
   "1101100001100000",
   "0001101000111100",
   "1110000011100011",
   "0010011000000100",
   "1101111111010110",
   "1110011011001100",
   "0010100010010010",
   "0010001001110000",
   "1101110011111101",
   "0010001111000011",
   "0001010101010111",
   "1101101111010101",
   "1101100100100000",
   "1101101001101101",
   "1110011010110011",
   "0010100100101110",
   "1110100001011111",
   "1110001001100000",
   "0010100101011001",
   "0010100100101011");



