
GS2 i LUTs

constant lut_gs : vector_of_std_logic_vector16(0 to 4095) := 
  ("0000000010001011",
   "0000000001110111",
   "0000000001000011",
   "1111111111110110",
   "1111111110011100",
   "1111111101001000",
   "1111111100001101",
   "1111111011111100",
   "1111111110101011",
   "1111111111110001",
   "0000000001000011",
   "0000000010010100",
   "0000000011010011",
   "0000000011110011",
   "0000000011101010",
   "0000000010110100",
   "0000000011100000",
   "0000000001010000",
   "1111111110010101",
   "1111111011001100",
   "1111111000011011",
   "1111110110101001",
   "1111110110010110",
   "1111110111111010",
   "1111111001001100",
   "1111111110100101",
   "0000000101011101",
   "0000001100110010",
   "0000010011001101",
   "0000010111010000",
   "0000010111100011",
   "0000010011000001",
   "0000000110111011",
   "1111111000000010",
   "1111100101001010",
   "1111001111101001",
   "1110111001001101",
   "1110100011101100",
   "1110010000111000",
   "1110000010001010",
   "1101111010100110",
   "1101110101101100",
   "1101110100111100",
   "1101110111010101",
   "1101111011100010",
   "1110000000000100",
   "1110000011100110",
   "1110000101000111",
   "1110000110001111",
   "1110000010010111",
   "1101111100000101",
   "1101110100100111",
   "1101101101100110",
   "1101101000111100",
   "1101101000100001",
   "1101101101111100",
   "1101111000001001",
   "1110001100001100",
   "1110100111110101",
   "1111001001111100",
   "1111110000101100",
   "0000011001101100",
   "0001000010010100",
   "0001100111111101",
   "0010001010011100",
   "0010100011010011",
   "0010110011011000",
   "0010111010010100",
   "0010111000100101",
   "0010101111001100",
   "0010011111100111",
   "0010001011011011",
   "0001110001111011",
   "0001011000111001",
   "0000111111000111",
   "0000100100110010",
   "0000001001101110",
   "1111101101100000",
   "1111001111110011",
   "1110110000101011",
   "1110001110100100",
   "1101101101100011",
   "1101010010010011",
   "1100111100111111",
   "1100110000001000",
   "1100101101111011",
   "1100110111111011",
   "1101001110101011",
   "1101110011101011",
   "1110011110001000",
   "1111010001001100",
   "0000000110001110",
   "0000111000001101",
   "0001100010010000",
   "0010000000001000",
   "0010001110110110",
   "0010001010110100",
   "0001110111001000",
   "0001011000100100",
   "0000110000011010",
   "0000000011001000",
   "1111010101101011",
   "1110101100111100",
   "1110001101010010",
   "1101110111110110",
   "1101110101010110",
   "1101111111111000",
   "1110011000110101",
   "1110111110000110",
   "1111101100011100",
   "0000011111111010",
   "0001010100001000",
   "0010000111000001",
   "0010110010000101",
   "0011001111101000",
   "0011011111111111",
   "0011100010011111",
   "0011010111100101",
   "0011000000101110",
   "0010100000001001",
   "0001110110010111",
   "0001001001000010",
   "0000011101110000",
   "1111110100111010",
   "1111010000101101",
   "1110110010110101",
   "1110011100100110",
   "1110001110111001",
   "1110001000001000",
   "1110001011001011",
   "1110011010011111",
   "1110110011001001",
   "1111010011110101",
   "1111111010101011",
   "0000100101010110",
   "0001010001001010",
   "0001111101010111",
   "0010100100010101",
   "0011000000101110",
   "0011010010101001",
   "0011011000110001",
   "0011010010101001",
   "0011000000101110",
   "0010100100010101",
   "0001111101010111",
   "0001010001001010",
   "0000100101010110",
   "1111111010101011",
   "1111010011110101",
   "1110110011001001",
   "1110011010011111",
   "1110001011001011",
   "1110000011110001",
   "1110001011001011",
   "1110011010011111",
   "1110110011001001",
   "1111010011110101",
   "1111111010101011",
   "0000100101010110",
   "0001010001001010",
   "0001111001000001",
   "0010100000100111",
   "0010111110101000",
   "0011010010111110",
   "0011011011111001",
   "0011011000011001",
   "0011001000010101",
   "0010101100011101",
   "0010001000101110",
   "0001011001000101",
   "0000100111011101",
   "1111110101011011",
   "1111000110111111",
   "1110100000000011",
   "1110000011111111",
   "1101110101010010",
   "1101110111011101",
   "1110000111101111",
   "1110100010000010",
   "1111000101111111",
   "1111110000001001",
   "0000011100100101",
   "0001000111010001",
   "0001101100100110",
   "0010001011111100",
   "0010100001000000",
   "0010101000110101",
   "0010100110110101",
   "0010011101011101",
   "0010001111111100",
   "0010000001110100",
   "0001110110010011",
   "0001101101101001",
   "0001101011101110",
   "0001110010111101",
   "0001111111011000",
   "0010001101111110",
   "0010011010111111",
   "0010100010100111",
   "0010100001100010",
   "0010010011010110",
   "0001111110000000",
   "0001011011111000",
   "0000110001101101",
   "0000000011001000",
   "1111010100011000",
   "1110101001101000",
   "1110000110011010",
   "1101101111010100",
   "1101100010101011",
   "1101011101011001",
   "1101100000000101",
   "1101101000010101",
   "1101110011010010",
   "1101111110001001",
   "1110000110100010",
   "1110001101000011",
   "1110001010011110",
   "1110000101101111",
   "1101111101111110",
   "1101110101001010",
   "1101101101101111",
   "1101101010001100",
   "1101101100101100",
   "1101111000111111",
   "1110001101000110",
   "1110100110010010",
   "1111000101110101",
   "1111101010010001",
   "0000010001101000",
   "0000111001101011",
   "0001100000000011",
   "0010000100110000",
   "0010100011001011",
   "0010110111001011",
   "0011000010001000",
   "0011000011110110",
   "0010111100101100",
   "0010101101011110",
   "0010010111010100",
   "0001111101110000",
   "0001011111100101",
   "0000111011110001",
   "0000010110001111",
   "1111110000110111",
   "1111001101011011",
   "1110101101100101",
   "1110010010101110",
   "1101111011101001",
   "1101101011011110",
   "1101100100110000",
   "1101100100011101",
   "1101101001001001",
   "1101110001000000",
   "1101111010000010",
   "1110000010011001",
   "1110001010110010",
   "1110001011100111",
   "1110001011001010",
   "1110000111100110",
   "1110000001111001",
   "1101111011011111",
   "1101110101111111",
   "1101110010110101",
   "1101110000110110",
   "1101110011000010",
   "1101111011011111",
   "1110000110100000",
   "1110010001110111",
   "1110011011000000",
   "1110011111100100",
   "1110011101110001",
   "1110010111000110",
   "1110001001100100",
   "1101110100100110",
   "1101011101110110",
   "1101001001101100",
   "1100111100110010",
   "1100111011001110",
   "1101000111111010",
   "1101100001101101",
   "1110001110001001",
   "1111000011011000",
   "1111111110011111",
   "0000111001000001",
   "0001101100000011",
   "0010010001001100",
   "0010100011100000",
   "0010100010011111",
   "0010000111101001",
   "0001011100100001",
   "0000100100100001",
   "1111100111001001",
   "1110101100110111",
   "1101111101111011",
   "1101100001000111",
   "1101011000100110",
   "1101101000001011",
   "1110010000001011",
   "1111001000110000",
   "0000001001101110",
   "0001001001100010",
   "0001111110101111",
   "0010100001011001",
   "0010101110011010",
   "0010011101011101",
   "0001110111001001",
   "0000111110110110",
   "1111111100111000",
   "1110111011000110",
   "1110000011010111",
   "1101011110001001",
   "1101001110111011",
   "1101011010011011",
   "1110000001010001",
   "1110111011011010",
   "0000000000000000",
   "0001000100100110",
   "0001111110101111",
   "0010100101100101",
   "0010110101011011",
   "0010100101100101",
   "0001111110101111",
   "0001000100100110",
   "0000000000000000",
   "1110111011011010",
   "1110000001010001",
   "1101011010011011",
   "1101001010100101",
   "1101011010011011",
   "1110000001010001",
   "1110111011011010",
   "0000000000000000",
   "0001000100100110",
   "0001111110101111",
   "0010100101100101",
   "0010110001000101",
   "0010100001110111",
   "0001111100101001",
   "0001000100111010",
   "0000000011001000",
   "1111000001001010",
   "1110001000110111",
   "1101100010100011",
   "1101010001100110",
   "1101011110100111",
   "1110000001010001",
   "1110110110011110",
   "1111110110010010",
   "0000110111010000",
   "0001101111110101",
   "0010010111110101",
   "0010101011110000",
   "0010100010100111",
   "0010000100001011",
   "0001010010110100",
   "0000010101101111",
   "1111010101101111",
   "1110011011111000",
   "1101110000001111",
   "1101010110100001",
   "1101011000010100",
   "1101101110110100",
   "1110011000111000",
   "1111010000101101",
   "0000001110110111",
   "0001001011100010",
   "0001111111100111",
   "0010100011100111",
   "0010110111010110",
   "0010111101001111",
   "0010110101010100",
   "0010100011101101",
   "0010001101100110",
   "0001111000011001",
   "0001101000110000",
   "0001100011111111",
   "0001101000100011",
   "0001110010111010",
   "0010000010100110",
   "0010010011101111",
   "0010100001111001",
   "0010101000110101",
   "0010100101001100",
   "0010010111010011",
   "0001111000011101",
   "0001010000111110",
   "0000100010000001",
   "1111110000001001",
   "1111000000100011",
   "1110011000010101",
   "1101111011111000",
   "1101110000011101",
   "1101110100110100",
   "1110000110000101",
   "1110100100101010",
   "1111001101100101",
   "1111111101000000",
   "0000101110110000",
   "0001011110101101",
   "0010000111000001",
   "0010100111100000",
   "0011000000110010",
   "0011001111011011",
   "0011010011000000",
   "0011001011101111",
   "0010111010100001",
   "0010100000101011",
   "0001111101110000",
   "0001011010011100",
   "0000110010010111",
   "0000001010000010",
   "1111100011101011",
   "1111000001001110",
   "1110100100001011",
   "1110001101100100",
   "1101111111111111",
   "1101111000100011",
   "1101110011111001",
   "1101110011001011",
   "1101110101001010",
   "1101111000100010",
   "1101111100000011",
   "1101111110100111",
   "1110000001101101",
   "1110000010010101",
   "1101111110001001",
   "1101111000001110",
   "1101110010000010",
   "1101101101011011",
   "1101101100010011",
   "1101110000011011",
   "1101111000111111",
   "1110001001011000",
   "1110100100001011",
   "1111000110001001",
   "1111101101011001",
   "0000010111011000",
   "0001000001010001",
   "0001101000001100",
   "0010000111011010",
   "0010100011101001",
   "0010110101000100",
   "0010111101100001",
   "0010111101010001",
   "0010110101000111",
   "0010100110001010",
   "0010010001101100",
   "0001111011000110",
   "0001100000110100",
   "0001000001001101",
   "0000011111100010",
   "1111111100111000",
   "1111011010011001",
   "1110111001010011",
   "1110011010110010",
   "1110000010010000",
   "1101101010000111",
   "1101011001110110",
   "1101001111110101",
   "1101001100011101",
   "1101001111110101",
   "1101011001110110",
   "1101101010000111",
   "1110000010010000",
   "1110011010110010",
   "1110111001010011",
   "1111011010011001",
   "1111111100111000",
   "0000011111100010",
   "0001000001001101",
   "0001100000110100",
   "0001111111011100",
   "0010010101011011",
   "0010101000010001",
   "0010110100110010",
   "0010111010001001",
   "0010110111110001",
   "0010101101011110",
   "0010011011100000",
   "0010000100110000",
   "0001100111101110",
   "0001000011010111",
   "0000011100000000",
   "1111110011111111",
   "1111001101101111",
   "1110101011011111",
   "1110001111000000",
   "1101110111010010",
   "1101101011011110",
   "1101100100110000",
   "1101100100011101",
   "1101101001001001",
   "1101110001000000",
   "1101111010000010",
   "1110000010011001",
   "1110000110011100",
   "1110000111111000",
   "1110001001000011",
   "1110000111111010",
   "1110000101000001",
   "1110000001010000",
   "1101111101100101",
   "1101111010111101",
   "1101110111110110",
   "1101110111001110",
   "1101111011011111",
   "1110000001100100",
   "1110001000001001",
   "1110001101101010",
   "1110010000101010",
   "1110010000000001",
   "1110001001000110",
   "1110000010110111",
   "1101110111111100",
   "1101101100011000",
   "1101100010100011",
   "1101011100110111",
   "1101011101011100",
   "1101100101110110",
   "1101111000111111",
   "1110010011111101",
   "1110110011000010",
   "1111010110101101",
   "1111111100111000",
   "0000100011001110",
   "0001000111011110",
   "0001100111101010",
   "0010000100010111",
   "0010010101111101",
   "0010100010100100",
   "0010101000000101",
   "0010100111001010",
   "0010100000111110",
   "0010010110111110",
   "0010001010111001",
   "0001111100001110",
   "0001101111001111",
   "0001100111110011",
   "0001100100011100",
   "0001100101010000",
   "0001101001111000",
   "0001110001100000",
   "0001111011000110",
   "0010000111100101",
   "0010001111000101",
   "0010010110111110",
   "0010011100000010",
   "0010011101011101",
   "0010011010101111",
   "0010010011101010",
   "0010001000001101",
   "0001111010101101",
   "0001100100101100",
   "0001001100111011",
   "0000110001011100",
   "0000010010100111",
   "1111110001000010",
   "1111001101101001",
   "1110101001110001",
   "1110001001010000",
   "1101100111011110",
   "1101001101000101",
   "1100111010000001",
   "1100110000001000",
   "1100110000111001",
   "1100111101001000",
   "1101010100110001",
   "1101111000111111",
   "1110100101000010",
   "1111010011010110",
   "0000000010101011",
   "0000101111010011",
   "0001010101100110",
   "0001110010010100",
   "0010000011000011",
   "0010001000100011",
   "0001111111111100",
   "0001100111101011",
   "0001000100011001",
   "0000011001100100",
   "1111101011010101",
   "1110111101111100",
   "1110010101010011",
   "1101110010010111",
   "1101011101110010",
   "1101010001101111",
   "1101001111111000",
   "1101010110100010",
   "1101100011000110",
   "1101110010011111",
   "1110000001101001",
   "1110001011110000",
   "1110010101101000",
   "1110010111111101",
   "1110010101010000",
   "1110001110101111",
   "1110000110001011",
   "1101111101100101",
   "1101110110110000",
   "1101110000110110",
   "1101101111000110",
   "1101110011111000",
   "1101111011110100",
   "1110000101000001",
   "1110001101010110",
   "1110010010110000",
   "1110010011101111",
   "1110001101011100",
   "1110000010110111",
   "1101110111111100",
   "1101101100011000",
   "1101100010100011",
   "1101011100110111",
   "1101011101011100",
   "1101100101110110",
   "1101110100101000",
   "1110010000001110",
   "1110110000111011",
   "1111010111000010",
   "0000000000000000",
   "0000101000111110",
   "0001001111000101",
   "0001101111110010",
   "0010000111000001",
   "0010010110011011",
   "0010100000011101",
   "0010100011011101",
   "0010100000100101",
   "0010011001011000",
   "0010001111101011",
   "0010000101010001",
   "0001111001100100",
   "0001110000011101",
   "0001101101010000",
   "0001101101101110",
   "0001110001010001",
   "0001110110110110",
   "0001111101001110",
   "0010000011001010",
   "0010000101100000",
   "0010000110010010",
   "0010000111110111",
   "0010001000000011",
   "0010000111000000",
   "0010000101000100",
   "0010000010101010",
   "0010000000001100",
   "0010000000001100",
   "0001111100010000",
   "0001111011000100",
   "0001111010011001",
   "0001111010001011",
   "0001111010011001",
   "0001111011000100",
   "0001111100010000",
   "0001111011110101",
   "0001111100011101",
   "0010000000100100",
   "0010000101011001",
   "0010001010001000",
   "0010001101110011",
   "0010001111011110",
   "0010001110011010",
   "0010001100100000",
   "0010000111010110",
   "0001111101001110",
   "0001110001111010",
   "0001100111100100",
   "0001100000011000",
   "0001011110010110",
   "0001100010101101",
   "0001101111111010",
   "0010000010010011",
   "0010010101000111",
   "0010100111100110",
   "0010110110010100",
   "0010111101110010",
   "0010111011000101",
   "0010101100010000",
   "0010001110100111",
   "0001101001111100",
   "0000111010100001",
   "0000000110110001",
   "1111010011110101",
   "1110100111000011",
   "1110000101010100",
   "1101110010011000",
   "1101101110001100",
   "1101111111100010",
   "1110011110000010",
   "1111001000010101",
   "1111111001011010",
   "0000101011011110",
   "0001011000100100",
   "0001111011010101",
   "0010010001110100",
   "0010010110111110",
   "0010000111101111",
   "0001101000000000",
   "0000111011010101",
   "0000000110100010",
   "1111001111000110",
   "1110011010011001",
   "1101101010111110",
   "1101001010111101",
   "1100110101110100",
   "1100101110001111",
   "1100110011010000",
   "1101000010110000",
   "1101011001111001",
   "1101110101101100",
   "1110010001001110",
   "1110110001001001",
   "1111001101101101",
   "1111101000111000",
   "0000000011001000",
   "0000011101001100",
   "0000110111110011",
   "0001010011010001",
   "0001101101000101",
   "0010001010110010",
   "0010100100000000",
   "0010111000101001",
   "0011000110001010",
   "0011001010001011",
   "0011000010111000",
   "0010101111011011",
   "0010010010011000",
   "0001100110110101",
   "0000110110010111",
   "0000000010110001",
   "1111010000101101",
   "1110100100111111",
   "1110000011111111",
   "1101110001000110",
   "1101110000011101",
   "1101111111100110",
   "1110011010011100",
   "1111000000001111",
   "1111101101000001",
   "0000011100010001",
   "0001001001011000",
   "0001110000010101",
   "0010001011111100",
   "0010011101010001",
   "0010100110101110",
   "0010100111001001",
   "0010100000100101",
   "0010010101101100",
   "0010001001011010",
   "0001111110011011",
   "0001110100101001",
   "0001101111111011",
   "0001110010111101",
   "0001111010011100",
   "0010000100010000",
   "0010001101101001",
   "0010010011101101",
   "0010010011110010",
   "0010001110000010",
   "0001111110110000",
   "0001100011011011",
   "0000111111100111",
   "0000010101101111",
   "1111101000111100",
   "1110111100101001",
   "1110010100000110",
   "1101110100001111",
   "1101011100010111",
   "1101001010111100",
   "1101000010011111",
   "1101000010101111",
   "1101001010111001",
   "1101011001110110",
   "1101101110010100",
   "1110001001010000",
   "1110100010111011",
   "1111000000111001",
   "1111100000001010",
   "0000000000000000",
   "0000011111110110",
   "0000111111000111",
   "0001011101000101",
   "0001111011000110",
   "0010010101011011",
   "0010101000010001",
   "0010110100110010",
   "0010111010001001",
   "0010110111110001",
   "0010101101011110",
   "0010011011100000",
   "0010000000011010",
   "0001100011111111",
   "0001000001010001",
   "0000011100010100",
   "1111110111000111",
   "1111010011011111",
   "1110110011000101",
   "1110010111001000",
   "1110000010101001",
   "1101110011011001",
   "1101100110110110",
   "1101011111001101",
   "1101011100010011",
   "1101011101111001",
   "1101100011100010",
   "1101101100100001",
   "1101111010000111",
   "1110000100011100",
   "1110010000100110",
   "1110011010110000",
   "1110100001010110",
   "1110100011001010",
   "1110011111100000",
   "1110010110011001",
   "1110000110011100",
   "1101110011111001",
   "1101100011100101",
   "1101010101110000",
   "1101001100110100",
   "1101001010111101",
   "1101010001101111",
   "1101100001111110",
   "1101111001011000",
   "1110011101011011",
   "1111000101100010",
   "1111110001000101",
   "0000011100101100",
   "0001000100101101",
   "0001100101100100",
   "0001111100001101",
   "0010001000100011",
   "0010000110110010",
   "0001110100011011",
   "0001010101010001",
   "0000101100001011",
   "1111111100111011",
   "1111001011110000",
   "1110011100111001",
   "1101110001111110",
   "1101010000100101",
   "1100111101001000",
   "1100110101110101",
   "1100111001110110",
   "1101000111010111",
   "1101011100000000",
   "1101110101001110",
   "1110001110100100",
   "1110101001000000",
   "1111000110000110",
   "1111100011001000",
   "0000000000000000",
   "0000011100111000",
   "0000111001111010",
   "0001010111000000",
   "0001110101110010",
   "0010001110100001",
   "0010100110000111",
   "0010111000010101",
   "0011000011000010",
   "0011000100011011",
   "0010111011010010",
   "0010100111010011",
   "0010001011011000",
   "0001100010101001",
   "0000110110010111",
   "0000000111101100",
   "1111011010011010",
   "1110110010010101",
   "1110010010111001",
   "1101111110110110",
   "1101111010000111",
   "1110000010100100",
   "1110010100111111",
   "1110110010000000",
   "1111010111010010",
   "0000000001111100",
   "0000101110110000",
   "0001011010100000",
   "0010000100010111",
   "0010100011000111",
   "0010111011010010",
   "0011001001010111",
   "0011001100110000",
   "0011000101101011",
   "0010110101000001",
   "0010011100010001",
   "0001111111011100",
   "0001011001111110",
   "0000110100011101",
   "0000001110101010",
   "1111101010010001",
   "1111001000110011",
   "1110101011011111",
   "1110010011001100",
   "1101111110010011",
   "1101110011100110",
   "1101101100010110",
   "1101101010001101",
   "1101101100010001",
   "1101110001010100",
   "1101110111111100",
   "1101111110101011",
   "1110000010000110",
   "1110000111111000",
   "1110001001000011",
   "1110000111111010",
   "1110000101000001",
   "1110000001010000",
   "1101111101100101",
   "1101111010111101",
   "1101111100001101",
   "1101111010111101",
   "1101111101100101",
   "1110000001010000",
   "1110000101000001",
   "1110000111111010",
   "1110001001000011",
   "1110000111111000",
   "1110000010000110",
   "1101111110101011",
   "1101110111111100",
   "1101110001010100",
   "1101101100010001",
   "1101101010001101",
   "1101101100010110",
   "1101110011100110",
   "1101111110010011",
   "1110010011001100",
   "1110101011011111",
   "1111001000110011",
   "1111101010010001",
   "0000001110101010",
   "0000110100011101",
   "0001011001111110",
   "0001111111011100",
   "0010011100010001",
   "0010110101000001",
   "0011000101101011",
   "0011001100110000",
   "0011001001010111",
   "0010111011010010",
   "0010100011000111",
   "0010000100010111",
   "0001011010100000",
   "0000101110110000",
   "0000000001111100",
   "1111010111010010",
   "1110110010000000",
   "1110010100111111",
   "1110000010100100",
   "1101111110011101",
   "1110000010100100",
   "1110010100111111",
   "1110110010000000",
   "1111010111010010",
   "0000000001111100",
   "0000101110110000",
   "0001011010100000",
   "0010000000000001",
   "0010011111011000",
   "0010111001001011",
   "0011001001101011",
   "0011001111111000",
   "0011001011011011",
   "0010111100100111",
   "0010100100011001",
   "0010000110011100",
   "0001011110001010",
   "0000110100011101",
   "0000001001101110",
   "1111100000100011",
   "1110111011011101",
   "1110011100100101",
   "1110000101011100",
   "1101111000111111",
   "1101110100010111",
   "1101110011111001",
   "1101111000000111",
   "1101111110111000",
   "1110000101111000",
   "1110001010111101",
   "1110001100010111",
   "1110000111000001",
   "1110000001100101",
   "1101110110100110",
   "1101101010010100",
   "1101011111011011",
   "1101011000110111",
   "1101011001010010",
   "1101100010101111",
   "1101111000011010",
   "1110010011011010",
   "1110111000101111",
   "1111100011011011",
   "0000001111110111",
   "0000111010000001",
   "0001011101111110",
   "0001111000010001",
   "0010001000100011",
   "0010001010101110",
   "0001111100000001",
   "0001011111111101",
   "0000111001000001",
   "0000001010100101",
   "1111011000100011",
   "1110100110111011",
   "1101111011101001",
   "1101010111010001",
   "1100111001110010",
   "1100100111010010",
   "1100100000111111",
   "1100100111010010",
   "1100111001110010",
   "1101010111010001",
   "1101111011101001",
   "1110100110111011",
   "1111011000100011",
   "0000001010100101",
   "0000111001000001",
   "0001011111111101",
   "0001111100000001",
   "0010001010101110",
   "0010001000100011",
   "0001111000010001",
   "0001011101111110",
   "0000111010000001",
   "0000001111110111",
   "1111100011011011",
   "1110111000101111",
   "1110010011011010",
   "1101110100000100",
   "1101011111000000",
   "1101010111001011",
   "1101011001001011",
   "1101100010100011",
   "1101110000000100",
   "1101111110001100",
   "1110001001101101",
   "1110010010010111",
   "1110010100010010",
   "1110001101000011",
   "1110000000101000",
   "1101110010000010",
   "1101100101000001",
   "1101011101011001",
   "1101011110011110",
   "1101101000010100",
   "1101111110010010",
   "1110100010000001",
   "1111001110100111",
   "0000000000000000",
   "0000110001011001",
   "0001011101111111",
   "0010000001101110",
   "0010011100000010",
   "0010100101010000",
   "0010100100101110",
   "0010011010101011",
   "0010001010110110",
   "0001111001100111",
   "0001101011010111",
   "0001100011100110",
   "0001100010010010",
   "0001101110011000",
   "0001111111101101",
   "0010010101001100",
   "0010101010010010",
   "0010111001111011",
   "0010111111010101",
   "0010110110111000",
   "0010100000111101",
   "0001110111011111",
   "0001000011111011",
   "0000001001000111",
   "1111001101100101",
   "1110011000100100",
   "1101110000111010",
   "1101011100000010",
   "1101011111001101",
   "1101110011111101",
   "1110011101111111",
   "1111010101011010",
   "0000010010100111",
   "0001001101000100",
   "0001111100100101",
   "0010011010011111",
   "0010100100110000",
   "0010010011101001",
   "0001101111110101",
   "0000111100001100",
   "0000000000000000",
   "1111000011110100",
   "1110010000001011",
   "1101101100010111",
   "1101011011010000",
   "1101100101100001",
   "1110000011011011",
   "1110110010111100",
   "1111101101011001",
   "0000101010100110",
   "0001100010000001",
   "0010001100000011",
   "0010100101001001",
   "0010100111101100",
   "0010010001001100",
   "0001100111001000",
   "0000101111010011",
   "1111110001001001",
   "1110110100011110",
   "1110000000011001",
   "1101011000000010",
   "1101000100111100",
   "1101000000101011",
   "1101001011000000",
   "1101011111011011",
   "1101111000001010",
   "1110001111001101",
   "1110011111011000",
   "1110100011000010",
   "1110011011101010",
   "1110001101000110",
   "1101111000011111",
   "1101100010100011",
   "1101010000110001",
   "1101001000010001",
   "1101001101000100",
   "1101100011011001",
   "1110001000010100",
   "1110110110100101",
   "1111101011111001",
   "0000100010011110",
   "0001010100000001",
   "0001111010101100",
   "0010010001110100",
   "0010010100011110",
   "0010000100111000",
   "0001100111011110",
   "0000111101110000",
   "0000001100110110",
   "1111011010100111",
   "1110101100111100",
   "1110001001000101",
   "1101110000110110",
   "1101101101001110",
   "1101111000010001",
   "1110010011000100",
   "1110111010111110",
   "1111101100001000",
   "0000100010000000",
   "0001010111110111",
   "0010001011011000",
   "0010110010000101",
   "0011001111101000",
   "0011011111111111",
   "0011100010011111",
   "0011010111100101",
   "0011000000101110",
   "0010100000001001",
   "0001110110010111",
   "0001001001000010",
   "0000011101110000",
   "1111110100111010",
   "1111010000101101",
   "1110110010110101",
   "1110011100100110",
   "1110001110111001",
   "1110001100011110",
   "1110001110111001",
   "1110011100100110",
   "1110110010110101",
   "1111010000101101",
   "1111110100111010",
   "0000011101110000",
   "0001001001000010",
   "0001110010000001",
   "0010011100011010",
   "0010111110101000",
   "0011010111111001",
   "0011100101100111",
   "0011100101110000",
   "0011010111001111",
   "0010111010001101",
   "0010001110000010",
   "0001011000010101",
   "0000011111111010",
   "1111100111100001",
   "1110110100011000",
   "1110001011011111",
   "1101110000111110",
   "1101100111100110",
   "1101110010100010",
   "1110001110000010",
   "1110110100011111",
   "1111100011100101",
   "0000010101101111",
   "0001000100111110",
   "0001101011100101",
   "0010000100110100",
   "0010001111101111",
   "0010001000100011",
   "0001101101101011",
   "0001000100101010",
   "0000010010100111",
   "1111011101110101",
   "1110101100111001",
   "1110000101111010",
   "1101101111111000",
   "1101100111001001",
   "1101110011000100",
   "1110010000000110",
   "1110111010111110",
   "1111101111000111",
   "0000100111001101",
   "0001011101111100",
   "0010001100010101",
   "0010110101010000",
   "0011001111101100",
   "0011011100110001",
   "0011011100101101",
   "0011010000101011",
   "0010111010100001",
   "0010011100011110",
   "0001111011000110",
   "0001010110000010",
   "0000101100110111",
   "0000000011111110",
   "1111011101011011",
   "1110111011001001",
   "1110011110101011",
   "1110001001001011",
   "1101111101010101",
   "1101110100010111",
   "1101110011111001",
   "1101111000000111",
   "1101111110111000",
   "1110000101111000",
   "1110001010111101",
   "1110001100010111",
   "1110001011010111",
   "1110000101010011",
   "1101111000101101",
   "1101101010000000",
   "1101011100010011",
   "1101010011000110",
   "1101010001101011",
   "1101011010100111",
   "1101110001011001",
   "1110001111001101",
   "1110111000101111",
   "1111101000010111",
   "0000011001100100",
   "0001000111010111",
   "0001101100111000",
   "0010000110000001",
   "0010010010001101",
   "0010001101101100",
   "0001110110100101",
   "0001010001101111",
   "0000100011010010",
   "1111110000010001",
   "1110111101111100",
   "1110010001000111",
   "1101101011010111",
   "1101010101101010",
   "1101001010001001",
   "1101001010001000",
   "1101010011011010",
   "1101100010110001",
   "1101110100100110",
   "1110000101010111",
   "1110010100011100",
   "1110011001010111",
   "1110011010000100",
   "1110010100111100",
   "1110001011100111",
   "1110000000011011",
   "1101110101111111",
   "1101101110101000",
   "1101101110001100",
   "1101101110101000",
   "1101110101111111",
   "1110000000011011",
   "1110001011100111",
   "1110010100111100",
   "1110011010000100",
   "1110011001010111",
   "1110010100011100",
   "1110000101010111",
   "1101110100100110",
   "1101100010110001",
   "1101010011011010",
   "1101001010001000",
   "1101001010001001",
   "1101010101101010",
   "1101101111101101",
   "1110010100110101",
   "1111000000000011",
   "1111101111111100",
   "0000100000001010",
   "0001001011111110",
   "0001101110111110",
   "0010000101100011",
   "0010001011001101",
   "0010000001110101",
   "0001101100111000",
   "0001001100010011",
   "0000100011010010",
   "1111110101101101",
   "1111000111101001",
   "1110011100111101",
   "1101111011000100",
   "1101011101100101",
   "1101001100001111",
   "1101000100111000",
   "1101000110100100",
   "1101001111101011",
   "1101011110000101",
   "1101101111011111",
   "1101111111011011",
   "1110001110011110",
   "1110011101011010",
   "1110101000011010",
   "1110101110001011",
   "1110101101110110",
   "1110100111000111",
   "1110011010010101",
   "1110000110011100",
   "1101101111111101",
   "1101011011111111",
   "1101001011000100",
   "1100111111111111",
   "1100111101010010",
   "1101000100111011",
   "1101010111111101",
   "1101110100000100",
   "1110011010011101",
   "1111001010111111",
   "1111111111010100",
   "0000110010011011",
   "0001011111000010",
   "0010000000001100",
   "0010010010000001",
   "0010010100011110",
   "0010000100101011",
   "0001100001111110",
   "0000110010101111",
   "1111111100111000",
   "1111000111001100",
   "1110011000100010",
   "1101110110111011",
   "1101100100100001",
   "1101100110000100",
   "1101111101101110",
   "1110100110001110",
   "1111011010011010",
   "0000010011110011",
   "0001001011100010",
   "0001111011011011",
   "0010011100100111",
   "0010101111001101",
   "0010110101101000",
   "0010101111100100",
   "0010100000100101",
   "0010001101010010",
   "0001111010100000",
   "0001101100011111",
   "0001101000010101",
   "0001101000100011",
   "0001110010111010",
   "0010000010100110",
   "0010010011101111",
   "0010100001111001",
   "0010101000110101",
   "0010100101001100",
   "0010010111010011",
   "0001111000011101",
   "0001010000111110",
   "0000100010000001",
   "1111110000001001",
   "1111000000100011",
   "1110011000010101",
   "1101111011111000",
   "1101101100000110",
   "1101110001000110",
   "1110000011111111",
   "1110100100111111",
   "1111010000101101",
   "0000000010110001",
   "0000110110010111",
   "0001100110110101",
   "0010010010011000",
   "0010101111011011",
   "0011000010111000",
   "0011001010001011",
   "0011000110001010",
   "0010111000101001",
   "0010100100000000",
   "0010001010110010",
   "0001110001011100",
   "0001010111000000",
   "0000111001111010",
   "0000011100111000",
   "0000000000000000",
   "1111100011001000",
   "1111000110000110",
   "1110101001000000",
   "1110001010001110",
   "1101110001011111",
   "1101011001111001",
   "1101000111101011",
   "1100111100111110",
   "1100111011100101",
   "1101000100101110",
   "1101011000101101",
   "1101111000111111",
   "1110100001000110",
   "1111001011110000",
   "1111110111111111",
   "0000100010011110",
   "0001000111111011",
   "0001100101100001",
   "0001111001000010",
   "0010000011001111",
   "0001111100111110",
   "0001101101000111",
   "0001010010100111",
   "0000101111010011",
   "0000000101101010",
   "1111011000100011",
   "1110101011000111",
   "1110000010101001",
   "1101011111011001",
   "1101000001011000",
   "1100101101000010",
   "1100100100000111",
   "1100100111100111",
   "1100110111101011",
   "1101010011100011",
   "1101110111010010",
   "1110100110111011",
   "1111011000100011",
   "0000001010100101",
   "0000111001000001",
   "0001011111111101",
   "0001111100000001",
   "0010001010101110",
   "0010001000100011",
   "0001111000010001",
   "0001011101111110",
   "0000111010000001",
   "0000001111110111",
   "1111100011011011",
   "1110111000101111",
   "1110010011011010",
   "1101110100000100",
   "1101011111000000",
   "1101010111001011",
   "1101011001001011",
   "1101100010100011",
   "1101110000000100",
   "1101111110001100",
   "1110001001101101",
   "1110001110000001",
   "1110010000100011",
   "1110001010111101",
   "1110000000111101",
   "1101110101001010",
   "1101101010110001",
   "1101100100111111",
   "1101100110100111",
   "1101101111010100",
   "1110000010011110",
   "1110100010000001",
   "1111001001101100",
   "1111110110010010",
   "0000100100000011",
   "0001001111000101",
   "0001110011111110",
   "0010010010011000",
   "0010100010010010",
   "0010101010001010",
   "0010101000111001",
   "0010100000100101",
   "0010010011111100",
   "0010000101111110",
   "0001111001011010",
   "0001101110001110",
   "0001101100010001",
   "0001101101010000",
   "0001110010101010",
   "0001111010111111",
   "0010000100001100",
   "0010001100001000",
   "0010010000111010",
   "0010010011100000",
   "0010001100111110",
   "0010000100100001",
   "0001111001100000",
   "0001101110001001",
   "0001100101000000",
   "0001100000011100",
   "0001100010001111",
   "0001101000111010",
   "0001110110011100",
   "0010001011011010",
   "0010100010001010",
   "0010110110010100",
   "0011000011001110",
   "0011000100110010",
   "0010111000000110",
   "0010011001111101",
   "0001101110001001",
   "0000111010100001",
   "0000000001110101",
   "1111001010000111",
   "1110011001101101",
   "1101110110011010",
   "1101100100101000",
   "1101100100100001",
   "1101111100100100",
   "1110100011011111",
   "1111010110100011",
   "0000001111001001",
   "0001000101110011",
   "0001110011001011",
   "0010010001001001",
   "0010011101110000",
   "0010010100110111",
   "0001110101010001",
   "0001000101011110",
   "0000001100000001",
   "1111010000110011",
   "1110011011111000",
   "1101110100011011",
   "1101100001110111",
   "1101100100001011",
   "1101111000100001",
   "1110011110010100",
   "1111010000101101",
   "0000001001011011",
   "0001000001110101",
   "0001110011110001",
   "0010011100100111",
   "0010110110111000",
   "0010111111010101",
   "0010111001111011",
   "0010101010010010",
   "0010010101001100",
   "0001111111101101",
   "0001101110011000",
   "0001100110101001",
   "0001100111010100",
   "0001101101011101",
   "0001111001010011",
   "0010000111101110",
   "0010010100111011",
   "0010011101000111",
   "0010011101001000",
   "0010010101000010",
   "0001111101100010",
   "0001011101111111",
   "0000110110010100",
   "0000001001101110",
   "1111011011111101",
   "1110110000111011",
   "1110001100000010",
   "1101101101101000",
   "1101011101101110",
   "1101010101110110",
   "1101010111000111",
   "1101011111011011",
   "1101101100000100",
   "1101111010000010",
   "1110000110100110",
   "1110001101011100",
   "1110010000000001",
   "1110010000101010",
   "1110001101101010",
   "1110001000001001",
   "1110000001100100",
   "1101111011011111",
   "1101110111001110",
   "1101110011100000",
   "1101110111001110",
   "1101111011011111",
   "1110000001100100",
   "1110001000001001",
   "1110001101101010",
   "1110010000101010",
   "1110010000000001",
   "1110001001000110",
   "1110000010110111",
   "1101110111111100",
   "1101101100011000",
   "1101100010100011",
   "1101011100110111",
   "1101011101011100",
   "1101100101110110",
   "1101110100101000",
   "1110010000001110",
   "1110110000111011",
   "1111010111000010",
   "0000000000000000",
   "0000101000111110",
   "0001001111000101",
   "0001101111110010",
   "0010000111000001",
   "0010010110011011",
   "0010100000011101",
   "0010100011011101",
   "0010100000100101",
   "0010011001011000",
   "0010001111101011",
   "0010000101010001",
   "0001111101111010",
   "0001110100001100",
   "0001101111010110",
   "0001101101011010",
   "0001101110001001",
   "0001110001000110",
   "0001110101100111",
   "0001111011000010",
   "0001111110011111",
   "0010000010000101",
   "0010000111110111",
   "0010001100111111",
   "0010010000101110",
   "0010010010011011",
   "0010010001100100",
   "0010001101111100",
   "0010000101100000",
   "0001111011100000",
   "0001110011100001",
   "0001101100011111",
   "0001100111100100",
   "0001100101110100",
   "0001101000000011",
   "0001101110100100",
   "0001110110111010",
   "0010000010110001",
   "0010010011000001",
   "0010100010111111",
   "0010101111101110",
   "0010110110001100",
   "0010110011110001",
   "0010100110101000",
   "0010001011111101",
   "0001101011001011",
   "0000111111111101",
   "0000010000000100",
   "1111011111110110",
   "1110110100000010",
   "1110010001000010",
   "1101111010011101",
   "1101110100110011",
   "1101111110001011",
   "1110010011001000",
   "1110110011101101",
   "1111011100101110",
   "0000001010010011",
   "0000111000010111",
   "0001100011000011",
   "0010001001010010",
   "0010100110001010",
   "0010110101110111",
   "0010111010110011",
   "0010110110010100",
   "0010101010100101",
   "0010011010010100",
   "0010001000011001",
   "0001111001100100",
   "0001101101010110",
   "0001100010100110",
   "0001011100100010",
   "0001011011100010",
   "0001011111100000",
   "0001100111110011",
   "0001110011011011",
   "0010000011001111",
   "0010010011000001",
   "0010011110100101",
   "0010100110101110",
   "0010101010010010",
   "0010101000011001",
   "0010100000011101",
   "0010010010001111",
   "0010000000000001",
   "0001100111101010",
   "0001000111011110",
   "0000100011001110",
   "1111111100111000",
   "1111010110101101",
   "1110110011000010",
   "1110010011111101",
   "1101111000111111",
   "1101100101110110",
   "1101011101011100",
   "1101011100110111",
   "1101100010100011",
   "1101101100011000",
   "1101110111111100",
   "1110000010110111",
   "1110001101011100",
   "1110010011101111",
   "1110010010110000",
   "1110001101010110",
   "1110000101000001",
   "1101111011110100",
   "1101110011111000",
   "1101101111000110",
   "1101101100100000",
   "1101110011000010",
   "1101111011011111",
   "1110000110100000",
   "1110010001110111",
   "1110011011000000",
   "1110011111100100",
   "1110011101110001",
   "1110010111000110",
   "1110001001100100",
   "1101110100100110",
   "1101011101110110",
   "1101001001101100",
   "1100111100110010",
   "1100111011001110",
   "1101000111111010",
   "1101100001101101",
   "1110001110001001",
   "1111000011011000",
   "1111111110011111",
   "0000111001000001",
   "0001101100000011",
   "0010010001001100",
   "0010100011100000",
   "0010100010011111",
   "0010000111101001",
   "0001011100100001",
   "0000100100100001",
   "1111100111001001",
   "1110101100110111",
   "1101111101111011",
   "1101100001000111",
   "1101011100111100",
   "1101101011111001",
   "1110010010010001",
   "1111001000011100",
   "0000000110100110",
   "0001000011110001",
   "0001110111001001",
   "0010011001010001",
   "0010100011000100",
   "0010010101100010",
   "0001110101000010",
   "0001000100000110",
   "0000001001101110",
   "1111001110001100",
   "1110011001111000",
   "1101110100000010",
   "1101011111100110",
   "1101100001100101",
   "1101111011110101",
   "1110101000010000",
   "1111100000100011",
   "0000011100111011",
   "0001010101001110",
   "0010000010000001",
   "0010011111110101",
   "0010100100101110",
   "0010010110101001",
   "0001110101010110",
   "0001000101000010",
   "0000001011011110",
   "1111001111000110",
   "1110010110001101",
   "1101100011111110",
   "1101000010110101",
   "1100101110001110",
   "1100101000011111",
   "1100110000001000",
   "1101000010011011",
   "1101011100000000",
   "1101111001011010",
   "1110010101100101",
   "1110110001001001",
   "1111001101101101",
   "1111101000111000",
   "0000000011001000",
   "0000011101001100",
   "0000110111110011",
   "0001010011010001",
   "0001110001011100",
   "0010001110100001",
   "0010100110000111",
   "0010111000010101",
   "0011000011000010",
   "0011000100011011",
   "0010111011010010",
   "0010100111010011",
   "0010000111000001",
   "0001011110111010",
   "0000110100010000",
   "0000001000000001",
   "1111011101100010",
   "1110111000000101",
   "1110011010011111",
   "1110000110111110",
   "1110000001000111",
   "1110000110110001",
   "1110010100111111",
   "1110101101000101",
   "1111001101100101",
   "1111110100100110",
   "0000011111110110",
   "0001001100110000",
   "0001110110010111",
   "0010011100011010",
   "0010111110101000",
   "0011010111111001",
   "0011100101100111",
   "0011100101110000",
   "0011010111001111",
   "0010111010001101",
   "0010010010011000",
   "0001011100000011",
   "0000100010000000",
   "1111100111001100",
   "1110110001010000",
   "1110000101101110",
   "1101101001010111",
   "1101011111011110",
   "1101100111001011",
   "1110000110000111",
   "1110110010011001",
   "1111101000110101",
   "0000100010100101",
   "0001011000000100",
   "0010000010000101",
   "0010011010101100",
   "0010011100000100",
   "0010001011111110",
   "0001100110001000",
   "0000110001110100",
   "1111110110010010",
   "1110111011111010",
   "1110001010111110",
   "1101101010011110",
   "1101011100111100",
   "1101100110101111",
   "1110001000110111",
   "1110111100001111",
   "1111111001011010",
   "0000110111100100",
   "0001101101101111",
   "0010010100000111",
   "0010100111011010",
   "0010100010100111",
   "0010000100001011",
   "0001010010110100",
   "0000010101101111",
   "1111010101101111",
   "1110011011111000",
   "1101110000001111",
   "1101010110100001",
   "1101011000010100",
   "1101101110110100",
   "1110011000111000",
   "1111010000101101",
   "0000001110110111",
   "0001001011100010",
   "0001111111100111",
   "0010100011100111",
   "0010110111010110",
   "0010111101001111",
   "0010110101010100",
   "0010100011101101",
   "0010001101100110",
   "0001111000011001",
   "0001101000110000",
   "0001011111101000",
   "0001100100110100",
   "0001110000110011",
   "0010000010111010",
   "0010010110110111",
   "0010100111101010",
   "0010110000011011",
   "0010101101010100",
   "0010011001111101",
   "0001111000111011",
   "0001001110111000",
   "0000011101011010",
   "1111101001100100",
   "1110111000111101",
   "1110010001000010",
   "1101110110010000",
   "1101101001011100",
   "1101110010010100",
   "1110001001011011",
   "1110101110010001",
   "1111011100101110",
   "0000001111101111",
   "0001000010000100",
   "0001101110111001",
   "0010010000010011",
   "0010100110101000",
   "0010110011110001",
   "0010110110001100",
   "0010101111101110",
   "0010100010111111",
   "0010010011000001",
   "0010000010110001",
   "0001110010100100",
   "0001101010110110",
   "0001100101111100",
   "0001100110001001",
   "0001101010101100",
   "0001110010001111",
   "0001111011000111",
   "0010000011101000",
   "0010001100100000",
   "0010010010001000",
   "0010010001100100",
   "0010001101011111",
   "0010000111000000",
   "0001111111101001",
   "0001111000111101",
   "0001110100010101",
   "0001110000011111",
   "0001110100010101",
   "0001111000111101",
   "0001111111101001",
   "0010000111000000",
   "0010001101011111",
   "0010010001100100",
   "0010010010001000",
   "0010010000110110",
   "0010000111010110",
   "0001111101001110",
   "0001110001111010",
   "0001100111100100",
   "0001100000011000",
   "0001011110010110",
   "0001100010101101",
   "0001101011100100",
   "0001111110100100",
   "0010010011000001",
   "0010100111111011",
   "0010111001011100",
   "0011000011100010",
   "0011000010101011",
   "0010110100011000",
   "0010011001111101",
   "0001110001110111",
   "0000111100101000",
   "0000000001100001",
   "1111000110111111",
   "1110010011111101",
   "1101101110110100",
   "1101011100100000",
   "1101011101100001",
   "1101111000010111",
   "1110100011011111",
   "1111011011011111",
   "0000011000110111",
   "0001010011001001",
   "0010000010000101",
   "0010011110111001",
   "0010100111011010",
   "0010010111110101",
   "0001101111110101",
   "0000110111010000",
   "1111110110010010",
   "1110110110011110",
   "1110000001010001",
   "1101011110100111",
   "1101010101111100",
   "1101100110010010",
   "1110001010111110",
   "1111000000110110",
   "0000000000000000",
   "0000111111001010",
   "0001110101000010",
   "0010011001101110",
   "0010101010000100",
   "0010100001011001",
   "0001111110101111",
   "0001001001100010",
   "0000001001101110",
   "1111001000110000",
   "1110010000001011",
   "1101101000001011",
   "1101010100010000",
   "1101011101011001",
   "1101111011110101",
   "1110101101001100",
   "1111101010010001",
   "0000101010010001",
   "0001100100001000",
   "0010001111110001",
   "0010100101001001",
   "0010100011111110",
   "0010001111000110",
   "0001100111011100",
   "0000110010011011",
   "1111110110111001",
   "1110111100000101",
   "1110001000100001",
   "1101100011011001",
   "1101001100110111",
   "1101000010110001",
   "1101000101110000",
   "1101010010100110",
   "1101100101000100",
   "1101111000101101",
   "1110001001100000",
   "1110010110101101",
   "1110011000001110",
   "1110010100101001",
   "1110001011010100",
   "1101111110111000",
   "1101110010101011",
   "1101101010001100",
   "1101101000100000",
   "1101110001111110",
   "1110000100111110",
   "1110011110101011",
   "1111000000000101",
   "1111100111001001",
   "0000010001010100",
   "0000111011110001",
   "0001100011110010",
   "0010000100110000",
   "0010011111011100",
   "0010110101000100",
   "0011000010011101",
   "0011000110111110",
   "0011000010011101",
   "0010110101000100",
   "0010011111011100",
   "0010000100110000",
   "0001100011110010",
   "0000111011110001",
   "0000010001010100",
   "1111100111001001",
   "1111000000000101",
   "1110011110101011",
   "1110000100111110",
   "1101110110010101",
   "1101101100001110",
   "1101101100010011",
   "1101110010010111",
   "1101111011110000",
   "1110000101100100",
   "1110001101000011",
   "1110010000000101",
   "1110001111101101",
   "1110000101010011",
   "1101111000101101",
   "1101101010000000",
   "1101011100010011",
   "1101010011000110",
   "1101010001101011",
   "1101011010100111",
   "1101110001011001",
   "1110001111001101",
   "1110111000101111",
   "1111101000010111",
   "0000011001100100",
   "0001000111010111",
   "0001101100111000",
   "0010000110000001",
   "0010010010001101",
   "0010001101101100",
   "0001110110100101",
   "0001010001101111",
   "0000100011010010",
   "1111110000010001",
   "1110111101111100",
   "1110010001000111",
   "1101101111101101",
   "1101011001011000",
   "1101001100001111",
   "1101001001110100",
   "1101010000010010",
   "1101011101000001",
   "1101101100111111",
   "1101111101001111",
   "1110001001000110",
   "1110010001011100",
   "1110010111111101",
   "1110011010001100",
   "1110011000011100",
   "1110010011100001",
   "1110001100011111",
   "1110000100100000",
   "1101111110110110",
   "1101110101110011",
   "1101110000100010",
   "1101101101010001",
   "1101101100001010",
   "1101101101010001",
   "1101110000100010",
   "1101110101110011",
   "1101111010100000",
   "1110000000110010",
   "1110001010011001",
   "1110010011110110",
   "1110011011100100",
   "1110011111111100",
   "1110011111100100",
   "1110011001100100",
   "1110001011110000",
   "1101111101101101",
   "1101101010111001",
   "1101011000011010",
   "1101001001101100",
   "1101000010001110",
   "1101000100111011",
   "1101010011110000",
   "1101110001011001",
   "1110010110000100",
   "1111000101011111",
   "1111111001001111",
   "0000101100001011",
   "0001011000111101",
   "0001111010101100",
   "0010001101101000",
   "0010010001110100",
   "0010000000011110",
   "0001100001111110",
   "0000110111101011",
   "0000000110100110",
   "1111010100100010",
   "1110100111011100",
   "1110000100101011",
   "1101101110001100",
   "1101101001000010",
   "1101111000010001",
   "1110011000000000",
   "1111000100101011",
   "1111111001011110",
   "0000110000111010",
   "0001100101100111",
   "0010010000101100",
   "0010110001010101",
   "0011001000000101",
   "0011010010000101",
   "0011001111111000",
   "0011000011000001",
   "0010101101101101",
   "0010010010011101",
   "0001110001011100",
   "0001001111010101",
   "0000110000001101",
   "0000010010100000",
   "1111110110010010",
   "1111011011001110",
   "1111000000111001",
   "1110100111000111",
   "1110010000010001",
   "1101110110011100",
   "1101100001011100",
   "1101010000101010",
   "1101000101110111",
   "1101000010110011",
   "1101001000110101",
   "1101011000101001",
   "1101101111111001",
   "1110010100000110",
   "1110111100101001",
   "1111101000111100",
   "0000010101101111",
   "0000111111100111",
   "0001100011011011",
   "0001111110110000",
   "0010010010011000",
   "0010010111100000",
   "0010010101110100",
   "0010001101010101",
   "0010000001001000",
   "0001110100101100",
   "0001101011010111",
   "0001100111110010",
   "0001101001010011",
   "0001110110100000",
   "0010000111010011",
   "0010011010111100",
   "0010101101011010",
   "0010111010010000",
   "0010111101001111",
   "0010110011001001",
   "0010011100100111",
   "0001110111011111",
   "0001000011111011",
   "0000001001000111",
   "1111001101100101",
   "1110011000100100",
   "1101110000111010",
   "1101011100000010",
   "1101011111001101",
   "1101110011111101",
   "1110011101111111",
   "1111010101011010",
   "0000010010100111",
   "0001001101000100",
   "0001111100100101",
   "0010011010011111",
   "0010100100110000",
   "0010010011101001",
   "0001101111110101",
   "0000111100001100",
   "0000000000000000",
   "1111000011110100",
   "1110010000001011",
   "1101101100010111",
   "1101011011010000",
   "1101100101100001",
   "1110000011011011",
   "1110110010111100",
   "1111101101011001",
   "0000101010100110",
   "0001100010000001",
   "0010001100000011",
   "0010100000110011",
   "0010100011111110",
   "0010001111000110",
   "0001100111011100",
   "0000110010011011",
   "1111110110111001",
   "1110111100000101",
   "1110001000100001",
   "1101011111000011",
   "1101001001001000",
   "1101000000101011",
   "1101000110000101",
   "1101010101101110",
   "1101101010110100",
   "1110000000010011",
   "1110010001101000",
   "1110011001010111",
   "1110011000101100",
   "1110010010100011",
   "1110000110101101",
   "1101111000010010",
   "1101101011000101",
   "1101100010111001",
   "1101100010111000",
   "1101101010111110",
   "1110000010011110",
   "1110100010000001",
   "1111001001101100",
   "1111110110010010",
   "0000100100000011",
   "0001001111000101",
   "0001110011111110",
   "0010010010011000",
   "0010100010010010",
   "0010101010001010",
   "0010101000111001",
   "0010100000100101",
   "0010010011111100",
   "0010000101111110",
   "0001111001011010",
   "0001101110001110",
   "0001101100010001",
   "0001101101010000",
   "0001110010101010",
   "0001111010111111",
   "0010000100001100",
   "0010001100001000",
   "0010010000111010",
   "0010010011100000",
   "0010001100111110",
   "0010000100100001",
   "0001111001100000",
   "0001101110001001",
   "0001100101000000",
   "0001100000011100",
   "0001100010001111",
   "0001101101010000",
   "0001111010001011",
   "0010001101100001",
   "0010100001110110",
   "0010110011001100",
   "0010111101011110",
   "0010111101001011",
   "0010101111111110",
   "0010010010111101",
   "0001101001111100",
   "0000111010100001",
   "0000000110110001",
   "1111010011110101",
   "1110100111000011",
   "1110000101010100",
   "1101110010011000",
   "1101110010100010",
   "1110000011010000",
   "1110100000001001",
   "1111001000000000",
   "1111110110010010",
   "0000100101101110",
   "0001010000111101",
   "0001110011001100",
   "0010001010110100",
   "0010010010110010",
   "0010000111101111",
   "0001101100111100",
   "0001000101000010",
   "0000010011111000",
   "1111011110000000",
   "1110101000001001",
   "1101110100101000",
   "1101001101111011",
   "1100110000011000",
   "1100100000000001",
   "1100011101100001",
   "1100101000011011",
   "1100111111010010",
   "1101011111110111",
   "1110000101010011",
   "1110110011010000",
   "1111100000001010",
   "0000001011011010",
   "0000110010011011",
   "0001010010111011",
   "0001101011000001",
   "0001111001001111",
   "0001111010100011",
   "0001110101010011",
   "0001100011011010",
   "0001001000001111",
   "0000100101100110",
   "1111111101110000",
   "1111010011010110",
   "1110101001001110",
   "1101111111111111",
   "1101011100111001",
   "1101000100101110",
   "1100110110101001",
   "1100110011010000",
   "1100111010010101",
   "1101001010111111",
   "1101100011101111",
   "1110000100111010",
   "1110101001110001",
   "1111001101101001",
   "1111110001000010",
   "0000010010100111",
   "0000110001011100",
   "0001001100111011",
   "0001100100101100",
   "0001111010101101",
   "0010001000001101",
   "0010010011101010",
   "0010011010101111",
   "0010011101011101",
   "0010011100000010",
   "0010010110111110",
   "0010001111000101",
   "0010000011001111",
   "0001110111010111",
   "0001101111011010",
   "0001101010001100",
   "0001101000011000",
   "0001101010001100",
   "0001101111011010",
   "0001110111010111",
   "0010000011001111",
   "0010001111000101",
   "0010010110111110",
   "0010011100000010",
   "0010011101011101",
   "0010011010101111",
   "0010010011101010",
   "0010001000001101",
   "0001111010101101",
   "0001100100101100",
   "0001001100111011",
   "0000110001011100",
   "0000010010100111",
   "1111110001000010",
   "1111001101101001",
   "1110101001110001",
   "1110001001010000",
   "1101100111011110",
   "1101001101000101",
   "1100111010000001",
   "1100110000001000",
   "1100110000111001",
   "1100111101001000",
   "1101010100110001",
   "1101110100101000",
   "1110100001010011",
   "1111010001010000",
   "0000000011000000",
   "0000110010011011",
   "0001011011010110",
   "0001111001111011",
   "0010001011001100",
   "0010001011001101",
   "0010000000011010",
   "0001100101100100",
   "0000111111110001",
   "0000010010111111",
   "1111100011101111",
   "1110110110101000",
   "1110001111101011",
   "1101110100000100",
   "1101100010101111",
   "1101011001010010",
   "1101011000110111",
   "1101011111011011",
   "1101101010010100",
   "1101110110100110",
   "1110000001100101",
   "1110001011010111",
   "1110010000000101",
   "1110001101000011",
   "1110000101100100",
   "1101111011110000",
   "1101110010010111",
   "1101101100010011",
   "1101101100001110",
   "1101110110010101",
   "1110000100111110",
   "1110011110101011",
   "1111000000000101",
   "1111100111001001",
   "0000010001010100",
   "0000111011110001",
   "0001100011110010",
   "0010000100110000",
   "0010011111011100",
   "0010110101000100",
   "0011000010011101",
   "0011000110111110",
   "0011000010011101",
   "0010110101000100",
   "0010011111011100",
   "0010000000011010",
   "0001100000000011",
   "0000111001101011",
   "0000010001101000",
   "1111101010010001",
   "1111000101110101",
   "1110100110010010",
   "1110001101000110",
   "1101111000111111",
   "1101101100101100",
   "1101101010001100",
   "1101101101101111",
   "1101110101001010",
   "1101111101111110",
   "1110000101101111",
   "1110001010011110",
   "1110001000101101",
   "1110000010110011",
   "1101111100000011",
   "1101110011100111",
   "1101101011011101",
   "1101100101110101",
   "1101100100111111",
   "1101101010110011",
   "1101110110010101",
   "1110001010100110",
   "1110101001101000",
   "1111001111011100",
   "1111111001011010",
   "0000100100010111",
   "0001001100111110",
   "0001110000010000",
   "0010001001101011",
   "0010011110100100",
   "0010101000000100",
   "0010101001001110",
   "0010100011101101",
   "0010011001101100",
   "0010001101100100",
   "0010000001100010",
   "0001111001100100",
   "0001110100001100",
   "0001101111010110",
   "0001101101011010",
   "0001101110001001",
   "0001110001000110",
   "0001110101100111",
   "0001111011000010",
   "0010000010110110",
   "0010000101110100",
   "0010001001111110",
   "0010001100101010",
   "0010001101100110",
   "0010001100101010",
   "0010001001111110",
   "0010000101110100",
   "0010000010110110",
   "0001111011000010",
   "0001110101100111",
   "0001110001000110",
   "0001101110001001",
   "0001101101011010",
   "0001101111010110",
   "0001110100001100",
   "0001111001100100",
   "0010000001100010",
   "0010001101100100",
   "0010011001101100",
   "0010100011101101",
   "0010101001001110",
   "0010101000000100",
   "0010011110100100",
   "0010001110000010",
   "0001110011111110",
   "0001001111000101",
   "0000100100000011",
   "1111110110010010",
   "1111001001101100",
   "1110100010000001",
   "1110000010011110",
   "1101101010111110",
   "1101100010111000",
   "1101100010111001",
   "1101101011000101",
   "1101111000010010",
   "1110000110101101",
   "1110010010100011",
   "1110011000101100",
   "1110010101000001",
   "1110001101111010",
   "1101111110001100",
   "1101101011001001",
   "1101011000110110",
   "1101001011110101",
   "1101001000010001",
   "1101010001010000",
   "1101100110000011",
   "1110001100101101",
   "1110111100000101",
   "1111110001111110",
   "0000101000101110",
   "0001011010000110",
   "0010000000001100",
   "0010010110001110",
   "0010010111001001",
   "0010001001000101",
   "0001100111011110",
   "0000111000110100",
   "0000000011001000",
   "1111001101010001",
   "1110011110000010",
   "1101111011010101",
   "1101101011100010",
   "1101101101111111",
   "1101111111110100",
   "1110100000111110",
   "1111001101100101",
   "0000000000101100",
   "0000110101000001",
   "0001100101100011",
   "0010010000010011",
   "0010101011110010",
   "0010111101001011",
   "0011000010011001",
   "0010111100111001",
   "0010101111001100",
   "0010011100011011",
   "0010000111111011",
   "0001110010100100",
   "0001100001011111",
   "0001011000111001",
   "0001010111000110",
   "0001011011100010",
   "0001100100111100",
   "0001110001100000",
   "0001111111010010",
   "0010001010001111",
   "0010010011011111",
   "0010011100011110",
   "0010100010000111",
   "0010100011101101",
   "0010100000110011",
   "0010011001001010",
   "0010001100100111",
   "0001111001000001",
   "0001100101001010",
   "0001001010110100",
   "0000101100110101",
   "0000001100000001",
   "1111101001011100",
   "1111000110010101",
   "1110100100001001",
   "1110000110100110",
   "1101101000101100",
   "1101010010100010",
   "1101000011010100",
   "1100111100001010",
   "1100111101111000",
   "1101001000110101",
   "1101011100110101",
   "1101110110111010",
   "1110011100001110",
   "1111000100001111",
   "1111101110101100",
   "0000011000110111",
   "0000111111111011",
   "0001100001010101",
   "0001111011000010",
   "0010001001101011",
   "0010010011110010",
   "0010010011101101",
   "0010001101101001",
   "0010000100010000",
   "0001111010011100",
   "0001110010111101",
   "0001101111111011",
   "0001110000010011",
   "0001111010101101",
   "0010000111010011",
   "0010010110000000",
   "0010100011101101",
   "0010101100111010",
   "0010101110010101",
   "0010100101011001",
   "0010010010111101",
   "0001110100100001",
   "0001001001011000",
   "0000010111010101",
   "1111100011010100",
   "1110110010111001",
   "1110001011100010",
   "1101110001110110",
   "1101100110110010",
   "1101101110001000",
   "1110001001011011",
   "1110110011001101",
   "1111100110011100",
   "0000011101000101",
   "0001010000111110",
   "0001111100101001",
   "0010011110010011",
   "0010101101010100",
   "0010110000011011",
   "0010100111101010",
   "0010010110110111",
   "0010000010111010",
   "0001110000110011",
   "0001100100110100",
   "0001011111101000",
   "0001101000110000",
   "0001111000011001",
   "0010001101100110",
   "0010100011101101",
   "0010110101010100",
   "0010111101001111",
   "0010110111010110",
   "0010011111010001",
   "0001111011111001",
   "0001001001011011",
   "0000001111001011",
   "1111010011110101",
   "1110011110101001",
   "1101110110011010",
   "1101100000011100",
   "1101011101100001",
   "1101110100011011",
   "1110011011111000",
   "1111010000110011",
   "0000001100000001",
   "0001000101011110",
   "0001110101010001",
   "0010010100110111",
   "0010011101110000",
   "0010010001001001",
   "0001110011001011",
   "0001000101110011",
   "0000001111001001",
   "1111010110100011",
   "1110100011011111",
   "1101111100100100",
   "1101101000111000",
   "1101101000010111",
   "1101111000100001",
   "1110011001011000",
   "1111000110111111",
   "1111111100000101",
   "0000110010111011",
   "0001100110000001",
   "0010001110100111",
   "0010110000001011",
   "0011000010101011",
   "0011001000011110",
   "0011000011001001",
   "0010110101010001",
   "0010100001111011",
   "0010001100010100",
   "0001110101001110",
   "0001100101101011",
   "0001011000111001",
   "0001010010001010",
   "0001010001110101",
   "0001010111100110",
   "0001100010100110",
   "0001110001100010",
   "0010000100111011",
   "0010010100001111",
   "0010100100000001",
   "0010110000000000",
   "0010110110010100",
   "0010110101011000",
   "0010101100001011",
   "0010011010010011",
   "0010000010010010",
   "0001100010100101",
   "0000111010011110",
   "0000001110111011",
   "1111100011010100",
   "1110111011010011",
   "1110011010011100",
   "1110000011110011",
   "1101111011110011",
   "1101111100111101",
   "1110001101101100",
   "1110101010011010",
   "1111010000101101",
   "1111111101010101",
   "0000101100101010",
   "0001011010111110",
   "0010000010101011",
   "0010100111100000",
   "0011000000110010",
   "0011001111011011",
   "0011010011000000",
   "0011001011101111",
   "0010111010100001",
   "0010100000101011",
   "0001111101110000",
   "0001011010011100",
   "0000110010010111",
   "0000001010000010",
   "1111100011101011",
   "1111000001001110",
   "1110100100001011",
   "1110001101100100",
   "1101111011101001",
   "1101110100110101",
   "1101110001110011",
   "1101110011100000",
   "1101111000010010",
   "1101111110010011",
   "1110000011101001",
   "1110000110101111",
   "1110000100010111",
   "1110000010110011",
   "1101111100000011",
   "1101110011100111",
   "1101101011011101",
   "1101100101110101",
   "1101100100111111",
   "1101101010110011",
   "1101110110010101",
   "1110001010100110",
   "1110101001101000",
   "1111001111011100",
   "1111111001011010",
   "0000100100010111",
   "0001001100111110",
   "0001110000010000",
   "0010001110000010",
   "0010100010010010",
   "0010101010001010",
   "0010101000111001",
   "0010100000100101",
   "0010010011111100",
   "0010000101111110",
   "0001111001011010",
   "0001110010100100",
   "0001101111111111",
   "0001101111010110",
   "0001110010010110",
   "0001110111110111",
   "0001111110011100",
   "0010000100100001",
   "0010001000110010",
   "0010001000001010",
   "0010000101000011",
   "0010000010011011",
   "0001111110110000",
   "0001111010111111",
   "0001111000000110",
   "0001110110111101",
   "0001111000001000",
   "0001111001100100",
   "0001111101100111",
   "0010000101111110",
   "0010001111000000",
   "0010010110110111",
   "0010011011100011",
   "0010011011010000",
   "0010010100100010",
   "0010000100010111",
   "0001101101010010",
   "0001010010011011",
   "0000110010100101",
   "0000001111001001",
   "1111101001110001",
   "1111000100001111",
   "1110100000011011",
   "1110000010010000",
   "1101101000101100",
   "1101010010100010",
   "1101000011010100",
   "1100111100001010",
   "1100111101111000",
   "1101001000110101",
   "1101011100110101",
   "1101111011010000",
   "1110011111111101",
   "1111000110010101",
   "1111101110011000",
   "0000010101101111",
   "0000111010001011",
   "0001011001101110",
   "0001110010111010",
   "0010000010101011",
   "0010001111100101",
   "0010010011101101",
   "0010010010100101",
   "0010001101111110",
   "0010000111110010",
   "0010000001110111",
   "0001111101101011",
   "0001111001111101",
   "0001111101101011",
   "0010000001110111",
   "0010000111110010",
   "0010001101111110",
   "0010010010100101",
   "0010010011101101",
   "0010001111100101",
   "0010000010101011",
   "0001110010111010",
   "0001011001101110",
   "0000111010001011",
   "0000010101101111",
   "1111101110011000",
   "1111000110010101",
   "1110011111111101",
   "1101111111100110",
   "1101100000100100",
   "1101001010111100",
   "1100111101100011",
   "1100111001000010",
   "1100111101100011",
   "1101001010111100",
   "1101100000100100",
   "1101111111100110",
   "1110011111111101",
   "1111000110010101",
   "1111101110011000",
   "0000010101101111",
   "0000111010001011",
   "0001011001101110",
   "0001110010111010",
   "0010000111000001",
   "0010010011010100",
   "0010010101110100",
   "0010010010010001",
   "0010001010110110",
   "0010000010000010",
   "0001111010010001",
   "0001110101100010",
   "0001110010111101",
   "0001111001011110",
   "0010000001110111",
   "0010001100101110",
   "0010010111101011",
   "0010011111111011",
   "0010100010100111",
   "0010011101010101",
   "0010010000101100",
   "0001111001100110",
   "0001010110011000",
   "0000101011101000",
   "1111111100111000",
   "1111001110010011",
   "1110100100001000",
   "1110000010000000",
   "1101101000010100",
   "1101011010110000",
   "1101011011010010",
   "1101100101010101",
   "1101110101001010",
   "1110000110011001",
   "1110010100101001",
   "1110011100011010",
   "1110011101101110",
   "1110010001101000",
   "1110000000010011",
   "1101101010110100",
   "1101010101101110",
   "1101000110000101",
   "1101000000101011",
   "1101001001001000",
   "1101100011011001",
   "1110001100001111",
   "1110111110001011",
   "1111110110100101",
   "0000101111010011",
   "0001100001101100",
   "0010000111011111",
   "0010011011110101",
   "0010011110001001",
   "0010001011100101",
   "0001100100001000",
   "0000101111001101",
   "1111110011111111",
   "1110111010100010",
   "1110001010101111",
   "1101101011001001",
   "1101011101111010",
   "1101101011001001",
   "1110001010101111",
   "1110111010100010",
   "1111110011111111",
   "0000101111001101",
   "0001100100001000",
   "0010001011100101",
   "0010011110001001",
   "0010011011110101",
   "0010000111011111",
   "0001100001101100",
   "0000101111010011",
   "1111110110100101",
   "1110111110001011",
   "1110001100001111",
   "1101100111101111",
   "1101001100110111",
   "1101000010110001",
   "1101000101110000",
   "1101010010100110",
   "1101100101000100",
   "1101111000101101",
   "1110001001100000",
   "1110010010010111",
   "1110010100011111",
   "1110010010100011",
   "1110001011101001",
   "1110000010000000",
   "1101111000011011",
   "1101110001110011",
   "1101110000101000",
   "1101111000111111",
   "1110001001001011",
   "1110011110101011",
   "1110111011001001",
   "1111011101011011",
   "0000000011111110",
   "0000101100110111",
   "0001010110000010",
   "0001111111011100",
   "0010100000001101",
   "0010111100100111",
   "0011010000010111",
   "0011011001100101",
   "0011010111000001",
   "0011001000000101",
   "0010101101001000",
   "0010000101010101",
   "0001011001110000",
   "0000100111001101",
   "1111110100000010",
   "1111000100101011",
   "1110011101011100",
   "1110000001111110",
   "1101110100111001",
   "1101110101001100",
   "1110000101001001",
   "1110100101010110",
   "1111001111111011",
   "0000000000000000",
   "0000110000000101",
   "0001011010101010",
   "0001111010110111",
   "0010001010110100",
   "0010001011000111",
   "0001111110000010",
   "0001100010100100",
   "0000111011010101",
   "0000001011111110",
   "1111011000110011",
   "1110100110010000",
   "1101111010101011",
   "1101010010111000",
   "1100110111111011",
   "1100101000111111",
   "1100100110011011",
   "1100101111101001",
   "1101000011011001",
   "1101011111110011",
   "1110000100111010",
   "1110101101101101",
   "1111010101001111",
   "1111111011101110",
   "0000011111011101",
   "0000111111000111",
   "0001011001101110",
   "0001101110101101",
   "0001111011101011",
   "0010000111011101",
   "0010001100000111",
   "0010001100110101",
   "0010001010110110",
   "0010000111011110",
   "0010000011111101",
   "0010000001011001",
   "0010000010101010",
   "0010000001011001",
   "0010000011111101",
   "0010000111011110",
   "0010001010110110",
   "0010001100110101",
   "0010001100000111",
   "0010000111011101",
   "0001111011101011",
   "0001101110101101",
   "0001011001101110",
   "0000111111000111",
   "0000011111011101",
   "1111111011101110",
   "1111010101001111",
   "1110101101101101",
   "1110000100111010",
   "1101011111110011",
   "1101000011011001",
   "1100101111101001",
   "1100100110011011",
   "1100101000111111",
   "1100110111111011",
   "1101010010111000",
   "1101110110010101",
   "1110100010100010",
   "1111010110101100",
   "0000001100010010",
   "0000111110011101",
   "0001101000010100",
   "0010000101101000",
   "0010010011010000",
   "0010010001110100",
   "0001111111000011",
   "0001011010101010",
   "0000101011001010",
   "1111110110010010",
   "1111000010100101",
   "1110010110011100",
   "1101110111011001",
   "1101101011100010",
   "1101110001111011",
   "1110000111011011",
   "1110101011101010",
   "1111011010011010",
   "0000001110010111",
   "0001000001110101",
   "0001101111100100",
   "0010010101100111",
   "0010101110110000",
   "0010110111101111",
   "0010110100001011",
   "0010100111001010",
   "0010010100110111",
   "0010000001110100",
   "0001110010000110",
   "0001100110101001",
   "0001100011100110",
   "0001101011010111",
   "0001111001100111",
   "0010001010110110",
   "0010011010101011",
   "0010100100101110",
   "0010100101010000",
   "0010011100000010",
   "0010000001101110",
   "0001011101111111",
   "0000110001011001",
   "0000000000000000",
   "1111001110100111",
   "1110100010000001",
   "1101111110010010",
   "1101100011111110",
   "1101011010110000",
   "1101011011010010",
   "1101100101010101",
   "1101110101001010",
   "1110000110011001",
   "1110010100101001",
   "1110011100011010",
   "1110011101101110",
   "1110010001101000",
   "1110000000010011",
   "1101101010110100",
   "1101010101101110",
   "1101000110000101",
   "1101000000101011",
   "1101001001001000",
   "1101100011011001",
   "1110001100001111",
   "1110111110001011",
   "1111110110100101",
   "0000101111010011",
   "0001100001101100",
   "0010000111011111",
   "0010011011110101",
   "0010011110001001",
   "0010001011100101",
   "0001100100001000",
   "0000101111001101",
   "1111110011111111",
   "1110111010100010",
   "1110001010101111",
   "1101101011001001",
   "1101011101111010",
   "1101101011001001",
   "1110001010101111",
   "1110111010100010",
   "1111110011111111",
   "0000101111001101",
   "0001100100001000",
   "0010001011100101",
   "0010100010011111",
   "0010011111100100",
   "0010001001100110",
   "0001100001010111",
   "0000101100001011",
   "1111110000110101",
   "1110110110100101",
   "1110000100000111",
   "1101011100011001",
   "1101000100111100",
   "1101000000101011",
   "1101001011000000",
   "1101011111011011",
   "1101111000001010",
   "1110001111001101",
   "1110011111011000",
   "1110100111011000",
   "1110011111011000",
   "1110001111001101",
   "1101111000001010",
   "1101011111011011",
   "1101001011000000",
   "1101000000101011",
   "1101000100111100",
   "1101011100011001",
   "1110000100000111",
   "1110110110100101",
   "1111110000110101",
   "0000101100001011",
   "0001100001010111",
   "0010001001100110",
   "0010011111100100",
   "0010011110001001",
   "0010000111110110",
   "0001100010000001",
   "0000101111100001",
   "1111110111000111",
   "1111000000010010",
   "1110010010010101",
   "1101110011010001",
   "1101101001010000",
   "1101110011000100",
   "1110001100110101",
   "1110110101010010",
   "1111100111001001",
   "0000011100000111",
   "0001001101100111",
   "0001110101101100",
   "0010010001110100",
   "0010011000011010",
   "0010001111000010",
   "0001110100100001",
   "0001001011101000",
   "0000011000011111",
   "1111100000000110",
   "1110100111101011",
   "1101110001111110",
   "1101000101110011",
   "1100101000110001",
   "1100011010010000",
   "1100011010011001",
   "1100101000000111",
   "1101000001011000",
   "1101100011100110",
   "1110001001101001",
   "1110110011010000",
   "1111100000001010",
   "0000001011011010",
   "0000110010011011",
   "0001010010111011",
   "0001101011000001",
   "0001111001001111",
   "0001111110111001",
   "0001111001000010",
   "0001100101100001",
   "0001000111111011",
   "0000100010011110",
   "1111110111111111",
   "1111001011110000",
   "1110100001000110",
   "1101111101010101",
   "1101011100011011",
   "1101000110110101",
   "1100111011010001",
   "1100111001110110",
   "1101000001111011",
   "1101010010010011",
   "1101101001010111",
   "1110000111100100",
   "1110101000100010",
   "1111001000001101",
   "1111100111101111",
   "0000000110100110",
   "0000100100011110",
   "0001000001001101",
   "0001011100100111",
   "0001111000011100",
   "0010001101010010",
   "0010100000101011",
   "0010101111000010",
   "0010110111000001",
   "0010110111011100",
   "0010101111100101",
   "0010011111001111",
   "0010000100110000",
   "0001100011111111",
   "0001000001010001",
   "0000011100010100",
   "1111110111000111",
   "1111010011011111",
   "1110110011000101",
   "1110010111001000",
   "1101111110010011",
   "1101101111101010",
   "1101100100110000",
   "1101011111100001",
   "1101011111011011",
   "1101100011101010",
   "1101101011001000",
   "1101110100101001",
   "1110000001001000",
   "1110001000101001",
   "1110010000100110",
   "1110010101110100",
   "1110010111101000",
   "1110010101110100",
   "1110010000100110",
   "1110001000101001",
   "1110000001001000",
   "1101110100101001",
   "1101101011001000",
   "1101100011101010",
   "1101011111011011",
   "1101011111100001",
   "1101100100110000",
   "1101101111101010",
   "1101111110010011",
   "1110010111001000",
   "1110110011000101",
   "1111010011011111",
   "1111110111000111",
   "0000011100010100",
   "0001000001010001",
   "0001100011111111",
   "0010000100110000",
   "0010011111001111",
   "0010101111100101",
   "0010110111011100",
   "0010110111000001",
   "0010101111000010",
   "0010100000101011",
   "0010001101010010",
   "0001110100000110",
   "0001011000111001",
   "0000111111000111",
   "0000100100110010",
   "0000001001101110",
   "1111101101100000",
   "1111001111110011",
   "1110110000101011",
   "1110001110100100",
   "1101101101100011",
   "1101010010010011",
   "1100111100111111",
   "1100110000001000",
   "1100101101111011",
   "1100110111111011",
   "1101001110101011",
   "1101101111010100",
   "1110011010011001",
   "1111001111000110",
   "0000000110100010",
   "0000111011010101",
   "0001101000000000",
   "0010000111101111",
   "0010010110111110",
   "0010010110001011",
   "0001111111000011",
   "0001011010101010",
   "0000101011001010",
   "1111110110010010",
   "1111000010100101",
   "1110010110011100",
   "1101110111011001",
   "1101101011100010",
   "1101110001111011",
   "1110000111011011",
   "1110101011101010",
   "1111011010011010",
   "0000001110010111",
   "0001000001110101",
   "0001101111100100",
   "0010010001010001",
   "0010101011000001",
   "0010110101101000",
   "0010110100011111",
   "0010101010010010",
   "0010011010101000",
   "0010001001011010",
   "0001111010001111",
   "0001101101101001",
   "0001100111110010",
   "0001101011010111",
   "0001110100101100",
   "0010000001001000",
   "0010001101010101",
   "0010010101110100",
   "0010010111100000",
   "0010001110000010",
   "0001111011000010",
   "0001100001010101",
   "0000111111111011",
   "0000011000110111",
   "1111101110101100",
   "1111000100001111",
   "1110011100001110",
   "1101111011010000",
   "1101100000100100",
   "1101001010111100",
   "1100111101100011",
   "1100111001000010",
   "1100111101100011",
   "1101001010111100",
   "1101100000100100",
   "1101111111100110",
   "1110011111111101",
   "1111000110010101",
   "1111101110011000",
   "0000010101101111",
   "0000111010001011",
   "0001011001101110",
   "0001110010111010",
   "0010000010101011",
   "0010001111100101",
   "0010010011101101",
   "0010010010100101",
   "0010001101111110",
   "0010000111110010",
   "0010000001110111",
   "0001111101101011",
   "0001111001111101",
   "0001111101101011",
   "0010000001110111",
   "0010000111110010",
   "0010001101111110",
   "0010010010100101",
   "0010010011101101",
   "0010001111100101",
   "0010000010101011",
   "0001110010111010",
   "0001011001101110",
   "0000111010001011",
   "0000010101101111",
   "1111101110011000",
   "1111000110010101",
   "1110011111111101",
   "1101111011010000",
   "1101011100110101",
   "1101001000110101",
   "1100111101111000",
   "1100111100001010",
   "1101000011010100",
   "1101010010100010",
   "1101101000101100",
   "1110000010010000",
   "1110100000011011",
   "1111000100001111",
   "1111101001110001",
   "0000001111001001",
   "0000110010100101",
   "0001010010011011",
   "0001101101010010",
   "0010000100010111",
   "0010010100100010",
   "0010011011010000",
   "0010011011100011",
   "0010010110110111",
   "0010001111000000",
   "0010000101111110",
   "0001111101100111",
   "0001111001100100",
   "0001111000001000",
   "0001110110111101",
   "0001111000000110",
   "0001111010111111",
   "0001111110110000",
   "0010000010011011",
   "0010000101000011",
   "0010001000001010",
   "0010001000110010",
   "0010000100100001",
   "0001111110011100",
   "0001110111110111",
   "0001110010010110",
   "0001101111010110",
   "0001101111111111",
   "0001110010100100",
   "0001111001011010",
   "0010000101111110",
   "0010010011111100",
   "0010100000100101",
   "0010101000111001",
   "0010101010001010",
   "0010100010010010",
   "0010010010011000",
   "0001110011111110",
   "0001001111000101",
   "0000100100000011",
   "1111110110010010",
   "1111001001101100",
   "1110100010000001",
   "1110000010011110",
   "1101101010111110",
   "1101100010111000",
   "1101100010111001",
   "1101101011000101",
   "1101111000010010",
   "1110000110101101",
   "1110010010100011",
   "1110011000101100",
   "1110010101000001",
   "1110001101111010",
   "1101111110001100",
   "1101101011001001",
   "1101011000110110",
   "1101001011110101",
   "1101001000010001",
   "1101010001010000",
   "1101100110000011",
   "1110001100101101",
   "1110111100000101",
   "1111110001111110",
   "0000101000101110",
   "0001011010000110",
   "0010000000001100",
   "0010010110001110",
   "0010010111001001",
   "0010001001000101",
   "0001100111011110",
   "0000111000110100",
   "0000000011001000",
   "1111001101010001",
   "1110011110000010",
   "1101111011010101",
   "1101101011100010",
   "1101101101111111",
   "1101111111110100",
   "1110100000111110",
   "1111001101100101",
   "0000000000101100",
   "0000110101000001",
   "0001100101100011",
   "0010001011111100",
   "0010101000000011",
   "0010111011000101",
   "0011000010101110",
   "0011000000000001",
   "0010110100111100",
   "0010100100000001",
   "0010010000000011",
   "0001111001100100",
   "0001100101101011",
   "0001011000111001",
   "0001010010001010",
   "0001010001110101",
   "0001010111100110",
   "0001100010100110",
   "0001110001100010",
   "0010000100111011",
   "0010010100001111",
   "0010100100000001",
   "0010110000000000",
   "0010110110010100",
   "0010110101011000",
   "0010101100001011",
   "0010011010010011",
   "0010000010010010",
   "0001100010100101",
   "0000111010011110",
   "0000001110111011",
   "1111100011010100",
   "1110111011010011",
   "1110011010011100",
   "1110000011110011",
   "1101111011110011",
   "1101111100111101",
   "1110001101101100",
   "1110101010011010",
   "1111010000101101",
   "1111111101010101",
   "0000101100101010",
   "0001011010111110",
   "0010000111000001",
   "0010101011001111",
   "0011000010111000",
   "0011001111000111",
   "0011001111111000",
   "0011000101111111",
   "0010110010111011",
   "0010011000100010",
   "0001110110110000",
   "0001010110001111",
   "0000110010010111",
   "0000001110111110",
   "1111101101011001",
   "1111001110100100",
   "1110110011000101",
   "1110011011010100",
   "1110000101010011",
   "1101110111110011",
   "1101101100010110",
   "1101100101010001",
   "1101100010100011",
   "1101100011111110",
   "1101101001000010",
   "1101110000111011",
   "1101111000011011",
   "1110000100111010",
   "1110001110100000",
   "1110010110001000",
   "1110011010110000",
   "1110011011100100",
   "1110011000001101",
   "1110010000110001",
   "1110001000001000",
   "1101111000110110",
   "1101101011001000",
   "1101011110101110",
   "1101010101101110",
   "1101010010001011",
   "1101010101110110",
   "1101100001111010",
   "1101111000111111",
   "1110010111111000",
   "1110111010101000",
   "1111100001011001",
   "0000001001101110",
   "0000110000111000",
   "0001010100010010",
   "0001110001101011",
   "0010000101010101",
   "0010010101001101",
   "0010011011000001",
   "0010011010001011",
   "0010010100100011",
   "0010001100011001",
   "0010000011111101",
   "0001111101001101",
   "0001111011101001",
   "0001111001010001",
   "0001111100010111",
   "0010000001101101",
   "0010000111101110",
   "0010001100100000",
   "0010001110001101",
   "0010001011001011",
   "0010000100010111",
   "0001110010011100",
   "0001011011110101",
   "0000111110110010",
   "0000011100010101",
   "1111110101111110",
   "1111001101101001",
   "1110100101100100",
   "1110000010010000",
   "1101011111010101",
   "1101000101011111",
   "1100110100010001",
   "1100101101000000",
   "1100110000100101",
   "1100111111001110",
   "1101011000100000",
   "1101111000111111",
   "1110100001010011",
   "1111010001010000",
   "0000000011000000",
   "0000110010011011",
   "0001011011010110",
   "0001111001111011",
   "0010001011001100",
   "0010001111100011",
   "0010000100001000",
   "0001100111101011",
   "0000111111011101",
   "0000001111110111",
   "1111011101111111",
   "1110101111000010",
   "1110000111100011",
   "1101101000101101",
   "1101011010110100",
   "1101010111001011",
   "1101011110000111",
   "1101101100010001",
   "1101111101011010",
   "1110001101000110",
   "1110010111011101",
   "1110010111101011",
   "1110010011100001",
   "1110000101100000",
   "1101110010101110",
   "1101011111011011",
   "1101010000011100",
   "1101001010011000",
   "1101010000110011",
   "1101100111101111",
   "1110001000010100",
   "1110110110100101",
   "1111101011111001",
   "0000100010011110",
   "0001010100000001",
   "0001111010101100",
   "0010010001110100",
   "0010011000110101",
   "0010001000100111",
   "0001101001100100",
   "0000111101011011",
   "0000001001101110",
   "1111010100110110",
   "1110100101010110",
   "1110000000111101",
   "1101101110001100",
   "1101101100110000",
   "1101111010011000",
   "1110010111101100",
   "1111000001100011",
   "1111110011101110",
   "0000101001010100",
   "0001011101011110",
   "0010001110000010",
   "0010110000110111",
   "0011001010001100",
   "0011010110101101",
   "0011010110011101",
   "0011001010100110",
   "0010110101000001",
   "0010011000000100",
   "0001111000011100",
   "0001010001110101",
   "0000101100110111",
   "0000001000111001",
   "1111100111001001",
   "1111001000011111",
   "1110101101100101",
   "1110010110111011",
   "1110000110111111",
   "1101110111010101",
   "1101101110011101",
   "1101101001111001",
   "1101101001001001",
   "1101101011100100",
   "1101110000010101",
   "1101110110100011",
   "1101111011000101",
   "1110000011101100",
   "1110001001000011",
   "1110001100110110",
   "1110001110101111",
   "1110001110100110",
   "1110001100011111",
   "1110001000101101",
   "1110000101110111",
   "1101111101111011",
   "1101111000001001",
   "1101110011000001",
   "1101101111010010",
   "1101101101100101",
   "1101101110011100",
   "1101110010000100",
   "1101111010100000",
   "1110000100100000",
   "1110001100011111",
   "1110010011100001",
   "1110011000011100",
   "1110011010001100",
   "1110010111111101",
   "1110010001011100",
   "1110000100110000",
   "1101111001100001",
   "1101101010111001",
   "1101011101010110",
   "1101010011011010",
   "1101001111100100",
   "1101010011110101",
   "1101100001100000",
   "1101110110101110",
   "1110010101010011",
   "1110111101111100",
   "1111101011010101",
   "0000011001100100",
   "0001000100011001",
   "0001100111101011",
   "0001111111111100",
   "0010001100111001",
   "0010000110110010",
   "0001110100011011",
   "0001010101010001",
   "0000101100001011",
   "1111111100111011",
   "1111001011110000",
   "1110011100111001",
   "1101110110010101",
   "1101010100010011",
   "1100111111001110",
   "1100110101100000",
   "1100110110101110",
   "1101000001100111",
   "1101010100011001",
   "1101101101000101",
   "1110001011111010",
   "1110101000100010",
   "1111001000001101",
   "1111100111101111",
   "0000000110100110",
   "0000100100011110",
   "0001000001001101",
   "0001011100100111",
   "0001110100000110",
   "0010001001100100",
   "0010011110100100",
   "0010101111010110",
   "0010111010001001",
   "0010111101001101",
   "0010110111001011",
   "0010100111010111",
   "0010001011110001",
   "0001101000001100",
   "0001000001010001",
   "0000010111011000",
   "1111101101011001",
   "1111000110001001",
   "1110100100001011",
   "1110001001011000",
   "1101110100101000",
   "1101101100101100",
   "1101101010001100",
   "1101101101101111",
   "1101110101001010",
   "1101111101111110",
   "1110000101101111",
   "1110001010011110",
   "1110001101000011",
   "1110000110100010",
   "1101111110001001",
   "1101110011010010",
   "1101101000010101",
   "1101100000000101",
   "1101011101011001",
   "1101100010101011",
   "1101101111010100",
   "1110000110011010",
   "1110101001101000",
   "1111010100011000",
   "0000000011001000",
   "0000110001101101",
   "0001011011111000",
   "0001111110000000",
   "0010010111101100",
   "0010100101010000",
   "0010100100101110",
   "0010011010101011",
   "0010001010110110",
   "0001111001100111",
   "0001101011010111",
   "0001100011100110",
   "0001100010010010",
   "0001101110011000",
   "0001111111101101",
   "0010010101001100",
   "0010101010010010",
   "0010111001111011",
   "0010111111010101",
   "0010110110111000",
   "0010011100100111",
   "0001110011110001",
   "0001000001110101",
   "0000001001011011",
   "1111010000101101",
   "1110011110010100",
   "1101111000100001",
   "1101100100001011",
   "1101100001110111",
   "1101110100011011",
   "1110011011111000",
   "1111010000110011",
   "0000001100000001",
   "0001000101011110",
   "0001110101010001",
   "0010010100110111",
   "0010100010000110",
   "0010010100110111",
   "0001110101010001",
   "0001000101011110",
   "0000001100000001",
   "1111010000110011",
   "1110011011111000",
   "1101110100011011",
   "1101100001110111",
   "1101100100001011",
   "1101111000100001",
   "1110011110010100",
   "1111010000101101",
   "0000001001011011",
   "0001000001110101",
   "0001110011110001",
   "0010011100100111",
   "0010110110111000",
   "0010111111010101",
   "0010111001111011",
   "0010101010010010",
   "0010010101001100",
   "0001111111101101",
   "0001101110011000",
   "0001100010010010",
   "0001100011100110",
   "0001101011010111",
   "0001111001100111",
   "0010001010110110",
   "0010011010101011",
   "0010100100101110",
   "0010100101010000",
   "0010011100000010",
   "0010000001101110",
   "0001011101111111",
   "0000110001011001",
   "0000000000000000",
   "1111001110100111",
   "1110100010000001",
   "1101111110010010",
   "1101100011111110",
   "1101011010110000",
   "1101011011010010",
   "1101100101010101",
   "1101110101001010",
   "1110000110011001",
   "1110010100101001",
   "1110011100011010",
   "1110011101101110",
   "1110010001101000",
   "1110000000010011",
   "1101101010110100",
   "1101010101101110",
   "1101000110000101",
   "1101000000101011",
   "1101001001001000",
   "1101100011011001",
   "1110001100001111",
   "1110111110001011",
   "1111110110100101",
   "0000101111010011",
   "0001100001101100",
   "0010000111011111",
   "0010011011110101",
   "0010011110001001",
   "0010001011100101",
   "0001100100001000",
   "0000101111001101",
   "1111110011111111",
   "1110111010100010",
   "1110001010101111",
   "1101101011001001",
   "1101011101111010",
   "1101101011001001",
   "1110001010101111",
   "1110111010100010",
   "1111110011111111",
   "0000101111001101",
   "0001100100001000",
   "0010001011100101",
   "0010100010011111",
   "0010011111100100",
   "0010001001100110",
   "0001100001010111",
   "0000101100001011",
   "1111110000110101",
   "1110110110100101",
   "1110000100000111",
   "1101100000101111",
   "1101001000101010",
   "1101000010110001",
   "1101001010101100",
   "1101011100010011",
   "1101110010011010",
   "1110000111100111",
   "1110010111010000",
   "1110100000011000",
   "1110011011001100",
   "1110001111001101",
   "1101111101000110",
   "1101101001001001",
   "1101011000010110",
   "1101001111100101",
   "1101010010101100",
   "1101100110000011",
   "1110000111000101",
   "1110110001001000",
   "1111100010100110",
   "0000010110011100",
   "0001000111000011",
   "0001101110111110",
   "0010001001110000",
   "0010010110100100",
   "0010001101101100",
   "0001110110100101",
   "0001010001101111",
   "0000100011010010",
   "1111110000010001",
   "1110111101111100",
   "1110010001000111",
   "1101101111101101",
   "1101011001011000",
   "1101001100001111",
   "1101001001110100",
   "1101010000010010",
   "1101011101000001",
   "1101101100111111",
   "1101111101001111",
   "1110001101011100",
   "1110010101001010",
   "1110011010000100",
   "1110011001110111",
   "1110010101010100",
   "1110001101110001",
   "1110000100111001",
   "1101111100011000",
   "1101110011100000",
   "1101101101111000",
   "1101101110011100",
   "1101110010100001",
   "1101111001000000",
   "1110000000010111",
   "1110000111000011",
   "1110001011101011",
   "1110001011001011",
   "1110000111111100",
   "1110000100111100",
   "1110000000101100",
   "1101111100001000",
   "1101111000010001",
   "1101110110000010",
   "1101110110000000",
   "1101110110001010",
   "1101111100110110",
   "1110000010110010",
   "1110001001001010",
   "1110001110101111",
   "1110010010010010",
   "1110010010110000",
   "1110001111100011",
   "1110000110011100",
   "1101111010101111",
   "1101110000010101",
   "1101100110101000",
   "1101011111011011",
   "1101011100100011",
   "1101011111100011",
   "1101101001100101",
   "1101111000111111",
   "1110010000001110",
   "1110110000111011",
   "1111010111000010",
   "0000000000000000",
   "0000101000111110",
   "0001001111000101",
   "0001101111110010",
   "0010000111000001",
   "0010010110011011",
   "0010100000011101",
   "0010100011011101",
   "0010100000100101",
   "0010011001011000",
   "0010001111101011",
   "0010000101010001",
   "0001111001100100",
   "0001110000011101",
   "0001101101010000",
   "0001101101101110",
   "0001110001010001",
   "0001110110110110",
   "0001111101001110",
   "0010000011001010",
   "0010000101100000",
   "0010000110010010",
   "0010000111110111",
   "0010001000000011",
   "0010000111000000",
   "0010000101000100",
   "0010000010101010",
   "0010000000001100",
   "0001111011110101",
   "0001111000100010",
   "0001111000111101",
   "0001111010101101",
   "0001111101010011",
   "0010000000001001",
   "0010000010101010",
   "0010000100011000",
   "0010000010110110",
   "0010000000101010",
   "0010000000100100",
   "0010000000011101",
   "0010000000011011",
   "0010000000011101",
   "0010000000100100",
   "0010000000101010",
   "0001111110100000",
   "0010000000101010",
   "0010000000100100",
   "0010000000011101",
   "0010000000011011",
   "0010000000011101",
   "0010000000100100",
   "0010000000101010",
   "0001111110100000",
   "0010000000101010",
   "0010000000100100",
   "0010000000011101",
   "0010000000011011",
   "0010000000011101",
   "0010000000100100",
   "0010000000101010",
   "0010000010110110",
   "0010000100011000",
   "0010000010101010",
   "0010000000001001",
   "0001111101010011",
   "0001111010101101",
   "0001111000111101",
   "0001111000100010",
   "0001111011110101",
   "0010000000001100",
   "0010000010101010",
   "0010000101000100",
   "0010000111000000",
   "0010001000000011",
   "0010000111110111",
   "0010000110010010",
   "0010000101100000",
   "0010000011001010",
   "0001111101001110",
   "0001110110110110",
   "0001110001010001",
   "0001101101101110",
   "0001101101010000",
   "0001110000011101",
   "0001111001100100",
   "0010000101010001",
   "0010001111101011",
   "0010011001011000",
   "0010100000100101",
   "0010100011011101",
   "0010100000011101",
   "0010010110011011",
   "0010000111000001",
   "0001101111110010",
   "0001001111000101",
   "0000101000111110",
   "0000000000000000",
   "1111010111000010",
   "1110110000111011",
   "1110010000001110",
   "1101110110110100",
   "1101100111101101",
   "1101011110011111",
   "1101011100101101",
   "1101100000111111",
   "1101101001100000",
   "1101110100001000",
   "1101111110110011");



